`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JNgwlIbp7nsVgY42mWPPDREjeTkRvVmq6cImXMnwabdkS5Tasq5r+X+lET4QLAWqUo5PIzKeymMm
eDGT3Uh7aQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KmhLxj8EHEOLo1zO5qehU7ubT877CKw/5FLL6CgHdR5DnViakTEut7hB2uKKyhy9TCQTjQJLiNck
vAzPejbV51gIi4TrhvW+FmARfccnrWDcdQ3NjIl/4y7WjpNBq+6W8jpmjUTzCA94B995kEkKBY4s
zoQ1T8uTb6KWfLT96H8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aUIPdVZH/XUnXSugmBFdTsOgfmQTf8WFZkka+WhWyR+6KcRAIF1RL3TaA8IxVbd+kgKgJ7Xe/aZs
KYwMUDdXzDNdQM2qjNv56zv/ZXArLpKznhHSGBkOkBJT7hgdXYQcfcUERikypwjk9HKhW9vRxNgP
lyA6dmwxCoPkZKR2hmEB9CGc4kHOmRYpZrglxgr8SgiIQCovY972BBWPJytVpVelv2SuMzx1J+sF
sbd5zoeewxTi5X6iMc/MADJpvtK6FaSVnEPW/d9BD8FhXD1B+XB96k9Zl5UfoGvU2vO6LVwmo1sM
wvq9kwqlSoPkYaSEWHte4E/4Pasg5cWBSqiMxA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YwD177lDyINODaxNS1zF9tP8s5u8SOhqmJysK0vhXApIbPgdsmSbWWunH195eGlJ7b6WTgBzS/yB
o43ZzK4W7ATh53nEHncGvtUoxzlRZlWgGBG5uSuh8HTtZtT3syer/+mLfS+GFM0Fafq35w+bxZEJ
a41K8FeA9rw6YGww1ro=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TdSeIm96C3p3yJEuyJcH4g3sdbUlXEcicmswtOZncE3XXR6U5F0qRaU3ccmluKnT+MSRKLRT1+JN
LJg0JGdXPdEAActX6GG1kZ+1jkCoNb2Egi3Z+zc7TVP7fM9Y6GCgUjKc6OrrICODKya8m38DThx2
zB62NdVPqT6QqN5uDNFvYgqLyGNPGqYP9SU5oGFQIfUsaLvmc2nyHmEoEXfHISmFZi0FU6GQSpHQ
SSvoaJmdykThQCSG0tAI0aTOIGVjXhqctbukHrqIFmG5R7Ht7m65iwUNgzc0nCMVgyLN95BC1x5w
HxA2QF6S1/oCVAXey3QcHA6yl2tYMNZXJjWq3A==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P6qxu3v2Dh5lKvwl7WFIkCTBJUyu4vpLCdo+Z702IGYzsVnbM/dCjjH/c+tyIMk7JfyR5f8DdGa9
aFwoQqldtPabDEhwtuNycrGtKVHCZR7UpxMxCAp5S8p35AykgNNjxlLjw34LbZ5JdqBLUaDeakyd
ksvD1SMyIC5C9+NnyFFDon4Ctd8Xfp98De+4pf1KK33OZPcppgda2gDq3uNGJVhNFdHQj8uqFRGi
j5p9h44HnGIrJDhPACACCIeEwB8qQt3BVHh4nJCo+/dd6nYxt93exE8Ys6imyHAEY79pkBD3YzFm
vZcIEUSd3YULQXZ11lAMTgSW4EE+Qx0DnfCHnw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 91216)
`protect data_block
1ABMSU5YAGNrAAAAAAAAADISj0kybV7EWAw4WNGABabI9uP+56CNbT3/rqaM5j9BL7Ou6FKhDZUG
58URxKpZNg0Vx1JyDFob+PJlLnfl7m5dz4Ab2I6IeTiB09lbT/PUcY9pTVtjUoEr0RWQnl4sQJXU
medr3I7x0lY4ZVgU9NacX1ahzp9bPcXbrC5giTJe1l6gxLne1RD5kMCn+plRRIBp1nYxuCe1/KkS
7jI+yMUB/EEzqRJghTCj+fhpTQVPWEh9kKxKQdO1ku6jGsNAMatT6TfOLyBqZvEICSbHfCu/pt/g
VkJPkjTDoPsYvPveabDPj+MY5+rYhCwv5Zxg1Gojgau1JJeexxoH1XIBmi74mAS0xLi926bP4tZu
msmKyHYVmJy0bQMcxSIhqdIFvfmn12I01eduAGXYnMmEx5rkYsfq4YGUbGcCatokd3LcmnroFn5+
sSKU+9Moalw7aLo7CdciCZdPWXyqtqltg78cMcUPLNTtY0M9MtJad0VoA/6DLVgo3tEmCjCABe+t
l5jj8rFiM0k1wIn4uipOiwfN9j5oIjSngQIhNNlZh09vZ9kGMIbxI5SLVoDW3hbP/nPPocIu48xG
dbS3yy4mZAIVQXL30rBgKd8wBT9Kq0YnJdpX/P/djzrU1jb64uFGI8DNx9IgYHndXHtgk6WWy1k8
FntGO3dMIh+tHEL2DZ7R8t8hnxMcwuv1SyNTSIxivA+3x+ch00GUk7Fe5Z/knxImNGWYuviPFVG3
AI9C/6/ADtxQ0sREwNPHOiEVlBha/Q8twhAKAmUmwgLs2MvIuFZt9/Q6uv0IKvUz1fGTXjBCuFeg
wm5U1CYBmAQshLCMt9td3b/zHoQjJ5shwf2lws3L+izorzcs9uRl+Pwp1pjq0FR+nG0ZRHTrOwuE
fjHuc8ypASnCCm3tzh0BcYkW0AzEfslGDwS7yNInvh7BYY3REnlDlTHbn3V1ZW7j37fQyqw4uYnW
oryT9/hYcDLDJvwc8ZOh+Cguac4j73+cHYlZdxKFUcLZ9bx+Q5RwQcBZzYphX6htWBex+sVEqOQE
m07JixAxQ/672yqYVpLQNkSCb3hVsH1n68eJ4/aJ8rBZygktcLlhR6F16iC55OKhEDg5/HD9Kjiv
XXqx8DgIEuMzfDiq/JGpCByh9GSp+6EzqMLDdd6iUm8GCLxnqYimmrRz2a3yomYtN29XNH5RiLXO
k1vVdanzOKpXlvNubXv4I44yuAcU+sedYWU32KT9iwX+6i619f1WI2pOzCAZVW1iK17LoRwxjUfR
LtPK6qg0BGoKChxAcfrRO30GJO4Z2w6NYJXRkZulpulL7SJoZvbE/AtZIdjpL8GlLXdM/axUhT08
C5u4e5vDUGL2sf4uqpkptzvvVURbPMWVQ2P61AQXgEt8bHvU5Rde/WZmGAv50RrNVw5RywYL+GF5
wLxjxPKe4ed2allcwkUcwHZPgaiRbYX30JgJ6NgKW35NfVky53GjX+Uv5s//o/cnmdS7jgTXwOIS
+yb7Fg1TAZ6KYnk62LdeaWxK0GtriFECEUHFhWhe1bk2xvDKGUHCrrSvovacIe06+XFGRF69RB59
aXDkhdJZwCJOxewmvnAIHrjsOLZrccwXUpc5zfvaiEQmE4En60uEo700vj7w2gudNZtobX0HM8d1
g4iXgtqlTFTua4JUu5tWO3gXI9yIq5A54vFHcF4Ztf4q5DN3N+kn1Q+5GjIeYGthutFzugP6k1tW
aqBlrmLVPvy+B2aD0Npj4QN8mb55ZkXx/TpkSUmpje/jjpUp2z3EI2abpcrT4DpuJwBs8KY9FZIj
Ufc7KkIfYsp+lM9LVBXqAcdUeZhuUyPx7saGMtyLBTifH7/513PL3+g2wxrto5as3dFsl3ktbOCV
Av4aGwO1R56MQPt+ld7CIuWjs0fIaRnqOAAj5Lq976xDbknE6xFGAe2wLQhM8roKn5Q8YMXY9Rvx
CWupFTjE7bhpNk1gUxIF/ejVm6+EoDmIiw27wmjlIesShDO5k0VpvCSbXI7Xg8MT1HVAFHejEAvn
3q35P9X5EBWZ2jbemMeF3Ir/rVdOKDfduEIM4y6V+eFcpiem/GXWSAtecLDqRPe7EjVn5rHZ+qT+
zmcnUmP/ZSG94UQWH6r26OcXW08882hQKumzkqRk3YE4/mWhezYJ56oyBk2QfGjAswgB4C1IOuPG
amTGlQPmgSSPnvjryjenbCK6IeA3ivO6lsk/HT/rKXSz8dFWGDz3r82wqms+E0DMsFhn6aQ1CwQH
Spcc6N/xaslWyY9IiW7LazqRCWDUSw2HYLA4yhEIo7y4RY3Xoqzn8ChhC1HvfcBmCJ4TV7raTlrk
htS7k/cNZl1Vz62nSzbNfTL+zQk3ORkp8zYhYM9wwnN2FYGupT+NotukSfZpKsygw5Eacc48w6/L
kwK75Tu4pnoZEpQDFLhJ5OHNNJAcWCmHh9B8otKv64TpKRZXuRWNJzt4b56JpIrWiDGRXEpZlS6W
0KNzaGdrB9oh3gCiwo0piwahxfUMsgDD4ja5naq+I7A2EJJsxOnJN2j+My9oVP58jB7fhumkoNyo
s3YYAKqjIeFEDwixgbMuyReJa5HADk8GDscskUiyt0/0CeDK3IWTPqe4h5sTFN3F3NWiK+0n9Hbr
PJDQw7gMyiHfXJInwBd92jEmS6fn2c1hpQp9eAdDC7v6I7tzOmq3qjx46+SIInRpbZlefdvxpEAw
CJebo7hdh5GPrn+7HzRKHEbsfn7Im/MQxnN0Lw9OHwWXfZeAb0ISMRd1Yggmvk+qeRJNNtVaxflR
M8fU0fs+ga0kp9icRUq5aSs9gd3IUS3RufuljKLnGbuhQ3Phbpm4pCqKwPNClUPOZf4niNHdtJQ7
fuGulvPGhSKfQEEZZUi0weH4ecCEvcfkfBPJjZ9QdYHcp42s0hqH6kjEJoW8qCO45gz/SGJ8Zabe
oWY2qh2x/i+DS2oAzoysoLD+5jGK2NLHUVfGb7Ny8xNkQmfsbYPjRa77rJ5pBbUAFtMqrh2qoGfD
BremUhvKkJdEVFm9S3q+oGbixuVhjdqznwXVYg/SbMXBbT44U0AvUlhTC8W8+qFR2HvBPQcvDv09
0Yow+JfeY7UW7LXc0E10iieB1DbRehQa6dhDzv21BsMFhfhjHDGzK3Zen3StjovSu05UeSu7ssZQ
tpk6g9R5RBa5Umaq4xpCMezbh0KcEpji905wrmu7KM3t2DcGx0m6uixlebBptjR7mhdBK3FitRCX
dAQRFkLOzUU0KWTcXY34wQewCyKBg//tEPHgPzmku7ekB6/OAnsGQw2HdvRqGXhvLm3yNsUzmxUv
s5igV6/8yVszzMNonYfb3njElE4Bt/U5kq8KoC1G9v+qa0vDU566bdBFk7TWPhILiFspqEAju5h7
xJWyAzTjCuFvsHpdhrHQfxCOds/g8nNF+i//zhR4aikdEZKy8r4FAP9o6g3b/9VOnN0AOSHFZTPw
IUb9l/ncCn7LJxsC7oqBBoVBfF0fTRH0bSjcX+LU9SPOzs9lNWg9pilUNGqdFowiNkwfB9MX7hCY
vaDLxqwfntvTk/v8n+hSG1Sn9+ceE69/q6bsnJIXXx9hbPoPDf89LkvOkEZMNvWdb33IvsKqz+lF
Z1cdypz2evHhrBzA8eYd8gjygU3Wdzc1O5fMrW2WvAnFnDJE+mGfIoKZr9TNf4iqx3+Hrdl44USV
tJzbfNfe/NXxZ1jtY50DnAX8OTF63gxtOKiE6E2g4AU25JIwp6fTOKt4MD6V0wJti2Abh+Yk0O63
iTob8Hzde7SzCfBECPKl7lK09XZ3ecb8X4RS6IQv3cGEiVDXHq16GEotrAc40pgZT08kn6PzxUBa
icqEdP7EN1/dI7dg4fOFkr8kpcvJIxiGsCQguU7dN/VxTmMmVJqpGyiTwQjn7sAuhbZHxENgiLlW
TmjkoAhkpdsiFnj2RlUGeDDRp166uhn+qpXI1GDNKjwkrlu6zXEcwO12jNsb8OWERpw6OsxxyKeK
nvzNqqKbrp0FYneRHXKLWM9a0QOsMBcbriMIe4EI5D+/8B0Sds7csH3sM+VkUs8kmiesNcvXRsMl
x8cKVoHAQN64R8yQqjQ8IrSyn5JZ5TtZGTPwlqrAoeGdlfbkXK65DWBNKmPQNErugOSU/tKrafKh
1RBtYMOFvzQ5Axo0jGP7PObyWlBhOGNo/pCQoX6sx3G0Ky6GHXzmMablHmu+OKIObPrzIEk7tn0E
SOySw8vnX/nlJdNc7009eGf+Oyck2mhD/FILBMxXlE2tVEWzuD9LpG1y1EZFsKURjhpGslobde+X
Ucjua4mBzQcEgJYfGyvwTCrMEe5xlHG1DErppGtmhbDGnVTACmzcntiSQrVVGSthNNQeCFcznk/I
3jOLTyVdTrcjhHBbv5SP6dlS46weL5quO3p4b7dgaM3s3HWJyV1yDdBxkeTlCd3CrspI2hBcd3JU
3LVLUIL/gmZFJP/OLSPJ8/SU3Gx+LQmpUJNiuziHntwjb454B1eaw1WG1ebupaKj01u+Q8CYrnMP
CLuAJI/IbKG3TcSRhlB7G2+yw0tcTUIy4uS6Zi6CO9ED7FwP0Lba8CTRNK6aSp8VlWhoOmZxoCXk
oMdPTMrKza71GrywnxkeAIzzgxr/tSW/5Hhs39CzMZDMh2eZpw7YiP553ycVu0+f2xxnC5d5TU2R
zUtuayweJpTdjIzMGcXTTOc6QBFmLAn+6XFR7uzR7aEEl1iWy1e7H0y2Fy/nyN3+LAOUfPMUxqKw
DPQitnFmXPSaDiF0reJ/hwqHp6heBujIIWE6Cmc8HXqBU+1ofc+Z8ePuNylMZsA+50KKyWp9D575
mvkcksEMBl6ituhA0jQp0rQ+bsCacLcXRPqJ8GjcGyO//TvcWizhHjl4obD/Qwc+tx4XRic02Ldg
Bf5hT4q8SRTSgJ9YrdjUu2PdLvBm+jU1/mUgnJYRan6d/ciP9LQW1eSMTaTKKNYu87argHsonbrb
Wb1i9WD0RSujJM+Zv0N8J5nBZLIf/hgXYZOcT9rHdCEmzK1Y+p4p6nUhMVnDP0KkEWZ8emGVlkhk
wYn/m3hpLxZxdAO/57QPOQmV8HPOyIqOtx4cgubt/tgypzrc0NDSnRQefBZUF5gFGZ9XpmkLXvsM
cJi7mpUNHzhpo4HgzcKbNwOwbb2vMwhGuHEJVqz/pQGOcSXn8FErH/SPJya6mZPv1kzSQf0zWT61
kYb8cKikp9e9xpM3pGnJxHKAEaT4kwNgk5FW8pJZQwm9tH8uhRLyD61WcW71SN23YRQUqwVpnr6f
qDrk7bd/wCjKLJz+gB6lh6D5uhUL12uqmEZKPsU+8UT+TuMLIBpL6F57vPAJvXvbb05T/ltV1vQ1
Xt48VVhF62iV9gc9wVOd03lGFYIe+qiN13TL3nNAViCiD2XQqRoS2UK1fF+rXfeyrX//May63APM
btjGmeb+C7ZYnXDDnBCQRBxpeZDaocXtriYZqyxw7xeYoVcpFd04c+poG8XCWdaNBdDTENyIcocQ
ZwPYZlvzqSymykY2QfCQ63YOe3cXVl/o3MgdubmOfFFFbqv1sjGhHFA60KEBxHK7CKcF7ZoiKh57
fQJwIVs8t6VPhRc/of4mdV/YkPxdE+xWMBHPVFX86Lr/J/nVNEQCigNl+r+ICDTpl3Eb+wVsmKQC
znMmDocu6Fd3T6d1UNa/wPwLzE5+BvEDlIPWdXV9CxUxHiDgnooxlENlX/5lw6Oc8XZpfU+RTQBs
njcB0U1DptQ7CIuMVm14WMSH76ktOR4lf+6JWK18ZMLrEQ+U77DUe6ju6Zj2x1duizKbiGTPfmvA
eZNKaETko/H7LZPZCWJYagA5ldrHcg8d4Yw/05V4eXqv3u0RxRVUSRrON7MXb37vThunSza7T7TP
Ns2hIEqZwIL3VmMJ2HgPgdmkfV2bpHZkuRtcRH1+sxBCDM5K1qpNgvDAG5/S6T3i4eSeU6vH11wK
8v3t5lKDbpMRPa/tR26qpL+eDQaCEBqNVC0FmIEs9MuLYAy6oYzSwGqLnQ0mbrThQ3JTBVFU81Nt
1ybz/K7xXaPgLqH8G08iMhDTKYPnIrZkvMhK3WOo+ktcnravd8Iaylee5gBj230BFxQvTDjHRhEy
l7S+MSJXSDsD/Mn/faonrAgT1nAfNa6IPWoGICNFKJByJ2SEpJcbM4QlW17wKu2nAz69rQOGNNno
42mXZLcZzTDXEk2IyClIsvtv1lFJWfdkW0pQYYKpJnS6CejY+6+K4lAGBS50l59c0bEosZrqXa29
mxXNhrIfakm55hXdqeQ+ZOrntiZw7Uh3NKfv8m5cqaWxwjKUUKcR4XnTTSsWys5liKcLWJzKgToQ
WVr/43OJfElCqcGfHpM0UsRbpyApKkdV8ufIQxc2vVWiU+xqfeLgp03oDziNCrmBIyD9ADTykm+7
+buKsjfZP9nqvfecOiJTdAWaQLbAU96Fwlp9bb2YoJQcZhgfszMCM/63FBC7E9RVN6Os5M6yeT0A
TPxoOoCigkiV9gFn6ZNIj6LGWvTWZSbg4MjWkJliH7CXPULHNr3bTmRVRocJ9eU8M+4RaWrwl06a
uFDuoknsa1Vgt1B3pj4ClL70e3eD03w0PrU/joLTA2kyPGRq/P3+aaWXFx+ratuDjfddcp7buSdU
gXMTLX4pehMdQKYyWuriWOK4fHfzI/9PRKcF+zXJQHGvFiWb4ye+CkCp/RJ1eF329LHBxS31zEak
mTZKgwEtBlDoqj+en2Y04qjiz8WCA3vUSeUqWk3Y17YFSZpUxm6AYNg3qHNhF8nLc4Z+MNucI+7Z
7ICflvZuTFYrfKZGBR5KU3ouLSCTFnYolR0F9fpl3mYCLd5TpyNXqQIHtTom43V/nHROSmYZnDbX
4lKj91pHZ5AvQY+dGgWUn6jwHMpA6cBHvQ83zJespuVN8220uzLKQpTf+xj+N7mT7iOz8hhGG3WE
wRkdT6wf3TqdlZcc4cGbeLSNTODeTyntp2DvnZ1hHJbFQy2zerT+4A2LseiJ+ipgkrw3DMcpMj3e
bnO0pHoqfjbMCo32bs28XFExug0qrkXXZ0mju1gV99hLlZHgvL5JR5mRcHOATHVLnsbiCifIbKE0
igs3IvPt110UJNy3GkU6q9yMyXvdZaH8XunIVCeSpi0RDaRGwfi7/x7oeGgoLn39xs3Yh/oVuJA0
0TwYNzRcON4/jVAe5eaONuJmQIOsYmBIAGeWAocKDHcXsgTeIQ30dPpDtR2s8FZCwH+tVmfG0W4d
xUv82JgO/GI3OUNcC4SYD0vBLKjaOZszfzklOPpR8Jm2a/KAeYZjvRgKtj3iIp/xZSM8INHq5iFN
1nfQEWBm8cw+nAG4JZ7VmHKDMCFk3eDnF6rThWCXoHe7oKomDqukmnH9TCX25ca/OKO1uIkZ3dl0
w8+FSXGF4GpwnbzOAUw2p/oIKGLZWtjqrh8YeTYJKVVGfeS4LhW7ZJ0D1JRxtZlsKS7zBksCR0tR
OgS3SrnxOFTW+JPr0pW83xjSoA50q9fL/4WjY07KTs5A8ORz+bhg8gJwfgxxQCQ5de0oG8UIML2o
zynGPuZFkOgYS8ves3nZc2njIc58PeYcoGZPzeAU3/q+vG7Afn9hjUaZRG8foUif82+Hhd7UBuvN
o3WjLdOyPH1DkY26V8CwiHx9pQv7KQ6xe1rn7Io7/WQIpndGjQ8Ul2K23jEDhq3TZHK5o8lbXAKa
MgH7hBTWChwSHP2MHZFaguC5jEigrRabXQfMEIljjVPq0llDUfnX/qH22x3ZuAR8VQkH5G5kaJrx
k7hpIzRHgwBb/9EiOT4ro0H3jWmDORp9ZBvgpCfEX4Frr7W0iZ0SVaoyhQAA5rBN69faGQYL18Md
2X1mnI2V7cB34c4+5Ybc7UCqo+Q0ast305+1zHUQdQgnzUY+yDjb4YzT5hDpSxzO+cV12XtECFhh
mYX6umPMn5vaB2mQpVDonLWJYRwpgQRQoKuTLQnLMUBE+dv7/1AmuXCPEDTmzh+bqINsYzohf2IY
+o9/01xbC7HzjIwB091OQAFTp+giiyUFYPctsvR+WKUoJrFqzCsCKEkGH7cQKvJlPKN2PDyLgLX/
1eCR5v5kW0GhLDdk4enOB3kEmhE4rQHQEku8eFYJQ1A9//EYRvTNIh+J0wcZ4whN/vX+loerxVfn
h4cUWdzqEzkmi3XDqLM0cpxRkItr+ku+oMSS6JEBmNFhuUeS98D2jWwvuR01blI5aCpKC4A0YHem
pX8zAaEq7K392iqIEuqraX9yL5U3T5xeXe1o8XeAEcWdi+xVOAxTRdBMtALTdJV585Y8OpbUEPRL
N42vjt2C7CgIyFMsjhZkl5pXjvG8YyJI2uoJdeGl8Gsplp6KkB37DgZD+TIjPZlUsV7fVt7kYd2E
pjgyo3Q9lIbWsZTQOUP+Q9yDTszA7A1UhSiNppTGUfda0yoFTBM1ScFGFpVT8NE983d7Gq5PKuFb
q3QSfZmUmm+Z1pDOdueSctbwfmU963qD5AEsTvms1/PVSvSbatxSsUTSUsLw9DJVgnKs6YpPosFU
cJf9B95EHDk9vqtf4nvUPhD0dH7Ssrbf8XeHH9M6o1xbwSMdP5fNlJfx9y/J9fIqaqyQWIpOoJ62
uWtIZDnlWWwmrsEmvswnSI7U15fRY4aJm00frVFfHbibGyzOmkPjPan4gTHISXVrKpoionE2OO20
4C9Qpsm356yUlwmXr8LmZw+trhdaMEHcEkPHi8l2/Or8ilK8t0zKaWDIUguUem9qljaGwRJE1z5v
biaiJQWzTw269TnGWpme/oZF39bqm+toSmUOrxgq5b0HgMhvd8VPdh5a7xVtA9K+uZ4bxiUkQlWY
pBSILno9FxOHXVWUiIvhbjCPrh25fqrIMY+uMhutf54sG93IZXNEUkOYRcLGqAIz+Y17SJGaS8LQ
YQto7UrYeqOLckv/6GiorgvNb6l1dAWOPnwHmMJSMbKw1GC5iOhNsOiaifgqHqKtb1jinqrwAuS2
rKAtKBISN1WawdlgzRWWE4V+XnIs/n8c+DeVZ3GoAKbDrdTYrX3HCjlvvyf2tibAw3MlGHv3Pfze
i5mdbP/Fkkr/9Xj6pBbSL54GUPVALGxrpS449+5jWu5+TYA+t+aRCBpIQNBlJTCZS4YRMoVwa6hi
kSHD+AiP9FeBSZlhd0GdQIyzbFALdR7itacgPc1WrlSNInPU+JZcP37Iy3/YikUlBpDTu2PuO259
8B4ZEhxzLE7hAOxunDk4bbYT0MpoXlXKKtpJdHLQRS8bd0BynY/1qW4Rsxf1h5wHdTmp36Zwc7bH
N+pwMDWupscto5wNbkjBMkhLfLYy/K5umjgxDGmZ0fc/RWD+9Ntl+bloSdw5uAQg4xHHxwew8EdF
UrPRVqqct7t9Qg1aj2HCu63H99PwDso6N3wZgdBbL4pu+aWB6qHZeKC83opQX8VHVFVUUg7W+F4L
DLE4/VrWqa3mEdTv4evCdvAjFTrfKvk5NsRPA1L3F65MRVoScZaVD+ARh0vdm8MgCZTqnMo4W4LG
qGxnMVU5VZ38y55VINU2zcvCJbWcBZv/hbIP/uqbTN4qdMd9mBTSgTr3nRxpknWKkp0aNwAuZ3OT
3mBQg97HiC2PXmJS4/m4IaeC1wvQehkqJZjbQNX9zrYvI5IxyVbJV+bwpyzL2u/+qTjV7+6RXPNV
dYJCL3+AQetWiWZ4A6eKyDM96tspmEhFaqxSNouIgCRpEfcL4AhAVZ45WqYgyiWkvj8856b0ZIw+
uVi0fC+FT5ccBqF3NLdD3aZKyAR3R7HdUv1SAF1b1sHsbq2gpERFlkmXdom14XIRzCGMr1ftpfr5
ytF2PBaxDSL8eqtirPbHD90KPDX+mSbdvgPPvTg/txqmuZCUvbAqnaJDlSdH2MPql6qgHBlsGG3Q
ciPltKD/w5+Zaa/kHpS9AsA17A8BFiN15SB3XdjTlhfMhV/t0nP4dtqEpGjCNs9H8AgIdBDAYXuE
V7KjK00MKUOrSoswp85olI0XZZ7+Xx9aj749+Szp5oxplxTO7ic1DosrRQ6yhmzfMlCYqnV4xNmV
O+GB2AvCTNpp4D7b9vaquLG5MIeDtdHZsL/SgzxDDotraNXtkXC6FD0drSA07Sc8n/3TySxlaF/+
Lo/jrTP5BXr5qsAmyim8CQa81Gfz/KWLx8lyxxPPJFwYQXYpeBeRjeYGnSLRvPl5iEbeaOuaDwAj
xuo/LfGWsxtOBVh4ZZtn+vCsn+sztjYxeIApctbrgMkOQw6XoK+dGSOKezMF8mwZd1uJe9lStAAJ
6hu51lobxSTz8JneyoGjvlyOX0yjZn+mUDsF4j00idv8PDS3mo/To3vMi0GVwNJ393wmbTzMZOK5
wqNrxb+lbuoBYxnO8uJ+cPz3favYozfk/bXqmHODNwoJJoOjaukuyM7/KZN0jULhHhicB5rCHh3J
XE6cY0QQivwzogBbOGoOfU3kS6CCvqKUqQHVcl2iRlMkPhNd1fd4imYA7q36qlhLeo4Ve4g8aKOD
EqZq2P3Vqk2tZ796Qu/enblbXekenrFy/T+DhanHixdQIyn1HpkVvswNPNF8hRxzxAwviGxavK9u
c1T8IpPaq3w4LZVjAYu4j8QH39kk5BVsQKjYgtZcWaBbID84mZaCMdlwHjspy/ge4j8bEWDFafQc
lD7oVGhv7zlqXxnokwfkSaSocweeI6n5Oe6LhrRd5ohHtG04tQlVB58AiOr/KuXaoVNYA+ikRVLn
t8dLbsHiDrfjkhNNZ8M+XvFSweBNkKp19qYk8EbmKQ/3AaILpeb5XlcU8TMp1vFnFHjSSRDcIUKT
h3iRKhnxZfyzORoySV/mQ6Wb1xaGp0jLDm0f6Wsie4WUQ5i0HLR2yKQIxrPI1ATaMwACxT3g4Kts
1397FdQpKEE/I5f1u3gVOZEZvD5p5jnMH+E1FK/xq8da0V5slAYshzyZNL8xuzXSXpdvbE2v3TVE
ug4Hud1/T3Xkr3tp6WiCOuXoC5QNvzQVGUkEs1QsOi3TYIhiaK9H/uFNRr6RkNbMrK+hji39yqIW
vyc7o2EnWbDh4gK+PRJ8yZfSRHBT3BSyO+Ksa0oPike9/9eFPdXKbnKULnwQ4WSMrHIDZgGwiiRf
BcP4AZLshCHlpC4bP+m+CmGZr0aOu716WBXKxz6V54NHzN0rU3WRtpssJI94T4qJm7hIS7szhVUq
+JKyoWLi8K5b/TNFmtlgZe+JBuo1gwQJFm447vXZKRiysuLdT5LZNcrvTYDx4VzzkG6aUlrAPOoS
jnL2/yydk8l7qmfXdVVSF0KcA3OV4wRXzFovCbNo3T2+RbtP0e4mU/r4YfnLck9NNgGPTHne+kLk
CxcgvhOtkyQ00lhN6z03n4xn0CNvKFpyuj+Zp0u7eb7VLotBGb7LXcahbZzz0PVGGOmXyIPU9ngQ
KNQnEPSZLzSOrbZAd4uKvDp+vJ0R/UwXT/eDezaXFqVslqthC1aH2c0w45bLkVmIDV6oK+s9oU2l
vjXbMIVIr9KTz45eIgOsPRzAkb5fwGLEYxBL+1Wqm+HoKVomnFWrCxTdFWMvz37XK4PVC4IEXv89
hCHfBPCseCo/1TDsTiZFRibzfN/iGT6ICaFLzX/BRhOXipYUoOsDRqFltvVe/GmBsk5ikf9IPNkx
mIO8kTDpupORJeWcL0vsj16HztMgER5ZrQ9ve9zS2vhM2tId0wwepltqCjqRs+Yq0CRioS12h/i+
mRuMBLMFFfm+qwWOAh+PW9T7jNCGrtdfPbdg6BRb8x2waT837lqJYnSsr2veWiBfYj13gVwIw2Vq
E2bTLSaN3WlBKuVsIeYtFhHM5KWL7gx/1oaz1QwRT1jrixwbxe1H655RaMEaSsdqq7AdJfGKCYVd
5usdBQK1+TckLKBzlvjUnwn1+IXXi3m2NOoihfIv+R55fYQzK6457DIj91MgmbdGz6jVf88psUM9
Uttdtger3ZSichm2qDRc++sRyaqK5StOTmy86Ueo3gHwckYNjkyK6HXAX6TKtj5wEw0HElrKaN1D
Ds03uJE+4840RwQsrYWFK8/uQe4Y9JL43UBO1dVl10wwRk/MgZXu0CmF6jVINwQkg8hcYqNklo+o
A2Cpy1Dyn2QQ5aSqn25pQFKfZdXTM3NRFdM7B28SoRnKwA3Z2u28F/mm4grHuK7wdCTzZjai1uYZ
T403E6AjEr/D+Za6ONM7euAZ2mapDaVx287dEsQmV/doqCNu4ur8n90SGcZqGUW0o0LUv6v2WQRp
hjeWIjEd8B+6PFSCkqKK9wA8UJFscyzLbQWZvAJPtnerr8h9CDRiLJgvawQBVRb44vr9I/nQShQD
hciCDsvj4A8GP/Ga5hCxvVyfqUEYD/MKYpY3cxyimA7nR6+9Nxqhuvs/jQuphqJT+0A90oeTorDS
9bfWdUT7lfvPIiG8HSImSObPcvrs/dSdP/P/Sn59HOWd0ylD++o0gADSuExVUG3UlgyMBfICpkrL
uv+n57hh4EVBooP4yI3ZW9TFYeqe8nGrHzJFDFSidv8cwB84A09j9BulM2zZ807ej2AdZc2jtueQ
Sx1NeoSSrKashjXSs3DzYX9/dCAkMRnmqjQ4rCZDIaUQ7FfWCJP7baLFOId+dUW+vYpmXm1pIIm8
BytqdMaSbaB3COIlkAQDTD8wVu3WNGipXk6YmXer0B6lfECdf/cfSft8mtG+XmK6KvpH5zZTPm4K
oUmHLdz6LPX6tJaQZTg0w8XdABTfCKZ08vy3Ba4s6eXV7oc4rfUmb1s/jTqr9p9H9z37mAGzdRDn
/Nt6mYTI6byCsPjzrdRvHnW6kSUTn+vVY61Zz3S1xCZSmQV61vADP0N36+vAdX53DiFzYg33eMTb
Mgd1m5bXhDA/8p67dTM6lfFujityxjGmQ+U++qFwcOnHNth99KCmu52/bBT8++N1rsvcNQYgWQ3S
7KvFb5/HGLJh7VxvF63zStuvlHQmBpnsWiXKeRI/iNNnwZ1i+izKLJK3GWxMLRahBWAHneT+5GKm
WP81el1CHhEurICOv/pHR3XLtzwx0172Lwp4ge0GbGwxRouwc92HQ5N2bX5uzqEx/rN9znCjQwD/
p7SFoy6/Llld+/OlBGTa9mQoNZKCDqgjASboUh5u0jP9qbp4JorcH64fKChj1m7/Ud7t8cvyXUvt
73yEb9NNLl2uEY+jJ3anvcJjX2phwLYEcxZ3gJZ7kYd70Hj20BhVp/LqbXGaXKf+4A+DkrN5cCSB
bnJcu6CTOmzS81kJNJY7DmC0sezDpo6LPIp1JlcZHhIvoE/LlM49sEtGOA4hVgPx7uM2EUhTB9v6
F5cIaeqCteXMagn6Od0vdMrr2Ay29VkS0xItUQfl5aXon2/Rcy3NWsH91z9uO6uOWuoMtmZwZ1CX
f/1IiqHQfEv63iYjiO/kdGEjLq0MAprorIIiRVJCI/o9WzBHrgLt2HH+TjHCLoHqF35HOoOcA4jX
/nAO4gSDg2giRgXAKY9MadsHi9FwMLX+yq9DYOnaww7xFL0xQCQWlj4Mct4HhfxIlYSV49o+nuiQ
KsCf4lezGrZ2rKdaXlj25gw7ZRgvJpJd7BoIkkxZta331ImlbfI83pFJc7eVxKs9Cg3DYI18Z420
YnIIk0+tnzPF8Oq4cq3IOqO4xT2DkHfWwZ+0/HjC5b3AzeOLst9rdVGg66NM9STpcQBmz3oWSx1/
yc1vNc0D0N0Lp01anBHsnXnpZBrV/OVCIVSKlC7FHagCS6FaxnmbWvgHVOCDIGWFPahrQttZkM5M
pA6QGv8C8jT5he3dvUgrPFA+Cwhgqcf9ZmxRYXNOpWUdBHse9wJOnoXcw/jqOy8JnOAbTRF5r/+X
7l25/hJT3+2jc2K2HJ7U5jkUZCQIJcijT1p2a/qUG8a94slLNm5FnG8lbPa0EPn1cfe9xClB+ddl
60b+8cS0P9zzw4SyX5JcRKZS19xOAJLt7xFLDBEfHi4naEEFb7MhDdEioOLOWg+d3WHfABZGxc7u
9YH0V2e4hxbgJs5i97fGBveXRp7ph+ETH43aiZ8Cy8Kwv9hUtZcrg3uJFHhGDZF7t3G0kBAxmGql
XcxA7VClIl54Mlsdg1q20Q5kyEunlLdCVp78SxV2q/QHSw8p7jzplRhI+/GpL+ZHQIeXB2OQXqxq
ndbXn5dIsEU3u2Z2s+9vF4A2P8H8AHB8BIPvHD0N1TQEa6pDbH9xR89l1WmiV1jb+BQMURZI1Inf
VeLeKHnrQVnkpYoXVhVh2K0V3FK0u5f6MfhpBURgkVWQy2w5NGQueI7hiTpG5qEI+ohcqqWkatZ4
Wps9/JW8bpLO5O7Xmpda9xiq/xoPHi7GRh6zheac3jp2fgLjlSYPJ57CjZAGLNC81Rt9bDG1PY3F
FatCLdzhRNDJBujVHUgDHGFzh+W/PJo2q5NmOgrQD4dkZLrIUgs759TcbVYpxAW5+6Y2wqROd1uN
JGMXOpRtuJni+0eNNdgfEpGBASTw9YJuSHihdnbdnhQt9TpFeSzaFmMtrJiF+yLHG4QTtCBHDAK5
cFeqlSd+xBPOHvzWA06B/j+z4FYMRYrErSXWfd90CjhG/E72EbXG7YQqljTkEqdmLYXZV27kqf0M
g8iz1em7KuWgOxTTH471h9bn5ipm8rNOyw0hxfiTeFhkzXINzXADvXUMy3Hi0GHgNDzFU8T5aJie
oWxe4pY+8jgMAsdwe5QC7efyTz8ec+ZNneJhVkWg1vX50en4+BPMcOOFCsakJhDQ8NO15AwOo85h
i0qthdWNuanQTwli72VaZZEq5LvWW74s1iAsamu6LxuSiJOuvttSCgsIWPf0Mz7b8X/kZSIUBXqN
mpZv73KWPUt/ZTatUrHNel6i5mBzOcBlndVemJX6M9P/edJADKJy8jk8bL/Ngw3C6apxHrJQDDRM
ksGdxa6bXWMKB3ITbYLP0/Qlv7xhloDWPiCJO25WN1u1w3C0uKQi6UsSuD48L4FEvyWchSMo21V1
1UNkvsJ8se+uN9AqQwZ85EiCyBx8TMYqO9DZJj28HnTbP01vmAQxS61+rWSwyazS+7M4Nx+HiX2I
Nd6cHo9qlbiKo2DRUpGYm5ntztsnrU3oisRzJeD6n4RsuMej/VB2Ry8gxnbBOUig7H9mnEuAAIE+
yXWayoZFtsdbrWOwKhi/XNs7sEw9RW/zGKk6wGecuGQARZTtq1NN+8QPjqSqVmKIZfou216Tu+BG
1S403vG++Mze2z+y3Upk9PQgcz4FBIxVGsKFXJVqayxua2lBAMCp4PlMJqnnU+72f7HU4GGSjZsu
GY52AWYHie7kzFiVJDZgRiiG9Wx1ux6gV8sdPrbZSgsTDOospiTWuU3kguc1ron+Dt5a7RD6F88y
BQQBB0sSFMmA3T4V+2BuNp5XFx/CsozGgV4KB2A2/OWna9E7/2mXLy05iKGwCvzYgEyA8M2t5Qyt
SqW1Dyl98yAkM6cqnAg5n6916NUi565Svs7+DHlq95QbG0KIV5HBYHwh9Mai1QjlGQ+8kStwqTI8
OZfTDfx0IsxzTxct3xTPeqIiQ4jaiXJwCDXz3WvDLDDpdCDjPDS0i/Gdv5O0uaUYC/LFMnV+iJtP
1a7LlyQ9Vtw6BTYvZ6tkQxeehAYkYtrabpvqMPp0XdRkVeeLgubR4z5KM5GhJ3pYLh85ZePxPk5W
p1RP3rp10XLPxymTUwU8XX582VEmYA7Jmy4B26ca3ITjOw8jxZFyAK+qdX+D9qwaSb5XhCYsLpzA
V3RVVR3puu+2im2GITZRWjn9uhlHjJtUf74qVl06gDOPXjc6za35pUAwvE2+Ag1EwjO2Ggh8sKZO
6JRxdv/t4WvVRUzlKIix6p9ONeD8EO+ykqzZ76ncS3dwqEBwiI3XrlxOAE3iY64n1GaoXrrfXwIK
VnaEvVMqjcp3GfeSfc8dqygIXpDW2+FIeJCKsL01dhPl40KorblJpX0srzqF9MQDSWmFCbwaHdx7
xUBu5JH/KE951mNvKlK7yXs0SSYxdd4qKYnVxDl3J5614VHOrzlq73B03Tps+Mxrywb5Q5gKUjKf
5/gwTysXdTUs4NuR0uOh1aT2LTVv2XYpXEQgTL+HkOV9vA/shKzLZBvEUXpWvqmOsoZJs4t9bfK+
9JQF/JXssIZamv0d/LnXyibke9JqhROGP3BWKrlv2GKe0fVEqtivqMZ3/W80xPqpia4xLn8qxxH0
hdfyHTpLRjsK3O5I6uK/cboYsrFjnEdmaKDEXec2CXiXwvTCiyidAj+R2XGuzc9Z6auWwvE/KTp8
+5FB4HcxbzeiOcA5KrVrMoxIMtRSbYh3+tKhYugW7DEXcrZmAVhC7HhMbWA+T7NOSfub+o2seIVD
TUVnbIcTzDPN7KM1UtAZrpwXASPfZl1ARcHWwDTNopg0fqZUAoGE3uvzEtdJqNC52hzSWE2ckqjh
PQnJEXwJO8r6d/oEiCQpIoBgBHM2z1zE64DSNSJ1IaFtsiMUFqNXO9YgEkgoVMIESHl7DtG/7AEw
tHJOiqf7KGAduEAB73VEHaWlvj/H/TrYg9yIL+wgeDB2fWBdVKPy2LID6znABGbUAt/tEudCnRGT
fNhr17OkvqFlmyHSIuVpYcaaJBkgoTDLS8swscdqux+h5fCwTzfT7WSFM0nMA9rQEsbXRkeA6mpO
wuiAaRjojdx2L60hilpRF56t6JFga5G/deOyviiMUUqDRAXg47a7VZSD6Hb9nOz3o/+cHeBKT76B
tA6FTMEI6IG/C3N8gP+v//vKSVbqCbRMqRL95F4Bg0MfN2loiXAX1KbP6M/P31E4T9YPqAoWTrcp
+svGa+tV0rYl+02KpUanOiZ710p0Y86GctPWYeLVQahGizh2fJtM3B+kcetX86d9NzIdozxoI30k
31W3awxZOb187cM0CpR5iFScEgVVChHZUDCEbBNG080Spk575hNllxIeqm7/PnC3JdR+VYmxufFO
Y2NpzQIGcvDOfhWX04+JKOj9zFnG9ZrvWiIqoxI7ZQqyxtbliF1IaqF+Qw9DvQkkan+V7plQSHYc
TX+mljmbLUYE97FUJJb5uFuPjj7vLWiDaCgwcYvMXCyFzXZtxQv1c8ng+m21kBXXfuvnZMiCMfVm
Km6tOH6giKHYzTrLwz6P0mrydGUpe479SxEJmbprflt7ptS4IviJB87har1yqxnO+ixHXXgdQnxE
VhrIBRN8B8r9c8v1GKsqouCa39HDHWbIBLD9sz3pI0/QFJa8szTZQsKLlxxoVYypILDC4u5GbzaJ
JBiFwqn8Po7yaIrl7fcZTHVK6lZ2EBaUFTE8OCbIVbFGxP9b8SzPT5B7NA9tFrXYmawzMwfCvIHC
1M52zXiaALwoxWx7ANb9sY5fjixBUxDrrp9fnEy75U3rWeJsHDuW4W+xq4VhU2fS74kNuTrVXAAd
QTlHK/32Vr4SKIkpAyzX/l//Abpb2e4Yq7c+pVbcH61qQnpTLErdiMjl2mDaJy0GJYBFUXEakgX2
2mpH/EUgzGZJYhXSyv2pYWrkObqhoeqNOJH/bukw92AZYNMalm4ZjbpbjJHtVt1LxIyoOETj/tNQ
p33C4hXKLfyK0jYQc3SLA6kduOBRuqypghIPzz9L3QbZnVRy1cyJzgHNH3qSJfRKE5+FVy8iY+rf
Ii3Z2nxyO3NeHBEZ+SYS9x72hxeBwOgm9zw49CZw+ZZpenlEr4oAXR65TmcOM/lcPfkowxnU3M0S
GGkpLXRsqpPcVPQRPeCx3NDJn91XfyO84KlxO4jyvWSzUaI81Vw7+qroSEIyUVtUnLnipaYzzZ5V
JztcNmu55SCvOrcjgMMtbVDr0aKdpSlrokl83+wxuq6igBF1oLRQ9ZORdtuK499PmNFbOtMCBaWA
x97Jrsziu6iXukGdsd1PNXsyAocBJp88ym1uzzxjFRFgMm+NQhrxRX+XOUbJufknxsoDpcy/hNC7
Y9bUglmetdSo4oBeIDsM7M0LFqLBSlclAP/UzFbzxyRvGiiVmfePy7sA8aEuFLyU9Z+oXo19l718
S/5/X1iTGUawP81NuMBxbI6Jquo6ULAA+Avky4BEpPiO3xITxy7yg7d+IZ236K/gXhRCBYqL7fs3
5rgOK4cFPD8aVqCxlFIagKU5HjGUKBotnanj706ACIezcDD2+K6q2Cr9JCUsiDHWNWNHOcbR5sJr
R8eFF3HUL26niloENUpXNcxglhClRvWZC++b/JFPnY3Tk7so7GpkNMdXoASWkO7dMfPDTMekwnCj
szioNvncPCObCiNgMtkJimB2awYtZpj0+2SzRznegN0SNnprwJ8fj8DXVVT9xsidlFJGKwrtEuRw
p4o+fA9txzlXGW3AfaLSt1xnavACY+4+G+cExsLpMkB8wTxZtve5GVers9pB23tZS4isBe9zr6nB
8uzEXPa7m819c7caeix6ykV6xoS6xzgeLgYfjsmHlK5wesExHDN/xzY7q5KEPRtMusxqHq3lbYti
ohM6JfA///jx2muuGkwQ4h3uaOCSwIkqp6gO0Lg+IgMm7SSRCSPF4klp7QGH05NgOOzZrGzgtc6/
oh5KrZa3YtC4/PXqLCmYVriAfzLBIOgAgPCTEn6J1ucpgxRs9xQitYdmQ4rd+LAyjIhuRWySIIXN
GDj7MgYB4k45AN/3VYlyqSAgs5ye7ZBUDrPMiGbdcJTXQRDG1C/6hsXqwnbF5mNpag18h2LWhgt9
GlurlyXda27TPJAo9Qw+80YjfG7WWAPVFCBd8Os1WijG/V6NKqLZ1Qc7H+88ViN7W1ZxQ7q1qXbV
3wK6MP9hpMBWCaDKIexMqUZkQMQ4Q4SxiBAdeD8pdbfch6+YqN7xpB5eWMTSvOGKMgHqT7VaIqeo
jm+Di+DWQiirWbd6A+wmSK51y0+uYvOdH80EETAxkvvMa1CVHo9DuWQeZmIci+qF43jAbp2nfPK5
W8x2/pQmlfqCDxKVPq9tf1yUS6kt7kazKybf4Of8y+6Z2/WDkBNbnQn1y/X+gzd1OqF4Uoqo7tRV
8gWm7V8CmZuD1WS70M4+9/I4hJ+h2u3SJlP/c8ShaVHi/EmGM+qDN4yaB/K1nJAGC7eHXQJXJ0WA
BW8wkcrPWC70lbuD1a6hEK33eeOkF+lVhj4fhy42Mjk8rIkwGO5TqbYdmBMI9Hy/h3hhc+kKqeTm
XHicDhqZAZiF5AKbaslrUVf07gzkA3R3TNVn8+iyqWbzIFLA1piG1Gr4EygWA3y0gMY/KqYRZcFJ
let/tLIe+CBvcgirrW6aK6PtAgpOc0r70fXuZ/Rq4QlW9cvUJd59lEKFwbn2xKTopwZYufxZCS1c
b4IHGnGGbgfqcgEZ21DtQuZIXIVrimpcDXhSxEAJA8yGLu8g18CNs05G3MS71bHdZAQ8KcyVtRM6
OSGwWyYBV3gQSgOw7XTBdzcGiJ2znBHcpDGmJlXB9udE171Zj1VOQTTbXv3ZEAnn8feZ5XF67wM5
ISAMa3YV8dHO5egQHOVh2ak1UAAy2t8D/IAGs1hGXDHstHGxTey9bKmx6mb/oZAVoX5gEtUaA82e
eNR8kpx6M78ru4K7stRnkoNhR5MqTKsaSRZSJugaU+CtgQ7D89kzhU2OhDoNDm51q98uqBogDj4+
xHZxMRla/ebVHUvHm20rLi2krhi4ryMw3s1ESNgEhTUOJvxhd4yz+hJZ3nFCtrWK281JlwVDvQ5G
OFb6PiokQAyMMdB2A3fWmFaraM+HGJQRKRUNCW5PUs2SG1CvBvlB+1IpJzhWLrheACFI1trBbhDy
W/Jhf9ZiXqq5XdoMPfvzawgATcZ6p9lWinOkRA9H7N/FGTomZVPBMaZpDA6+1WKDg6Ub9y27I6Ia
GFKczUdwW2+2KDi647DyK9hfsXvBauju2Vp4KvAcxfKTglfnRc1RJSTlMQjHqi//tWonWCDLXO1Y
czT2XN7Ff3mkYYUUWIeH3NPApVrwcXuc7AcBcJ80KzHJBYKylnuy7F/qDaEynnBJYhlFxBAK+oFp
ndjSh5nMcTqRGRKySDu0sCFjj1xBoIu8vopcLewDT43RePUYQmoSZGldkLIc8E7FBp4phVgytxO+
cqaDy63UWIQ8U9RA6pNhpbBXxuCoi8EV3geUMKiJd/1+CGQBYdi7JGhvcHylOqw/8VF97f1YB/P3
2k6fzc04BY9Zrb80ToJstxyr928bfOAmean9m29D560umxAP5hsosxwW0M4XSnsC+I7yN1b9zsH1
BI+qo1lnuljwBloayh+v1+7O6M0WvKwNtHbKnwp46OKD0D+oDSzkab+2FTRcHMbepwZr3jX4XWZg
86OYzjuEH+H5eT3pd7jV+e4e54vsugnnOyTs4N/3yI/342JwVCQnkkx8mVoUW9HHjt6QN6CBY+ta
83I6GTWemE+ISgTVgk3kBtChLeTiUrSCEx8VfB3bnl1z0Q0/FlsUF4BjwEpnUlG99ydh7qk07DVV
xDMMelyU7JYwKaQCrLeWb9kFxd3pa/I4pXcONlL3z7bjPnIo/yVauXwzml/dkWDafor+SHbEDwcH
yUVPWD1UMNotEKaiEAwiBHDAA1tfiRGN9tsYaMHT0TR2/3i+ZEJp7CfTpb1kxVCEZ+qTzCPKERTJ
hSV3zGDPVsBtK3JU2yqXbN6mLWMG7kEXDYXvJWoJ5JGjsaf2ZpdhcDuUBwB4iJ2uNxJhizZWXDro
Oy46Y1QQvb4K7DUESUXT8liszGQm0lxGL7B32087wfvDBww4QkIZzPMcMh+iGdxKIaoXkfIVbqcu
cJTUKCswvWgZTeXhqp4I33P85Tfr8G8eXPC9+9Z/FEvv9TLSr60mb6mfuEWoJNjZaji1TL3Iv7Tn
3ScZxAs6DQe47Qxmtg/5sWH9fF2ZTnZ/Hc/l+Jx/VLfRbg0iw56TXlHifUPuYQQqkeyfEiq8P6mu
QjAoO76gSRId4RmQzZyVRl9F2riteili7PEHeRdaH/FV7spMiNNfr8cQMAtmhpCM4SrEPnDILmem
wJtl9R9uZLHnGZVslS4hhxQp/rKZ4RvdQ+SOrtWQlMH2x7c4Ho4zeQ4NMgReaXwhYvVGzgKg2NmC
IjVvAv9/BGEkNDCW6uOc7s8Gz6tgvBskq+3jcykmszgOZxbz7X3mKOOQn/OoB6/dFVUVjrjEhs+/
Jt9wnMaQOit/PgwNMEuixX38XCAtbias4XktBV4NNIsMSM3o9S2wR+g50q2CWl2R/ygWrq1aHi3h
1XfLP9PbLtgvigLag6sgPqyxLvfavldwnSdB9wqVHowUhxZ6QcFk7LLR75Q2vCf/YIMjKK0HWc3U
JT5UQXJYXv6Yr5ZTWGI+aR/cPap0YRr5eIO8VY6nqn8kq91JsKceVZVZnc/EGejjQq+QjbIEW+Z6
FeHCd0PWefxSC9RoixrpnChPCLkseRfpkXj3yaAC6CxxxI8G5f79GhkPAeTKhCWAkySn6qj2BAcN
AEEeX5PFq0DoGNu5smi0cUSVK6O8wyyw9qfGnDvboAMwOgYJk8tF2J2LAuRQm7B8zrFvDFkqfoth
UDhyjgjbgMT9i7lspWhhES7rULweVj+bf7OVyencfLR3asWKRHEmFW8yTnjPIxDrM/Hv+zr/Uo16
CQwtcRypwWcjnvSge9wbP8K10QVE6WVsgnRFDCtgahZWa859Tp1fDTnGnGVzXOlSHs9NwohGpUaJ
q5BKKkzUQai1FOto2wfO2bftr+8w2vO8rdYjdCYXyznZN9idT/Jog3EDlatHC2FZSzwEzvOL/GL8
DQIlcrL1ZWdYt25Z3OMNSR8LftbttsGVcHqD9MiUrJSQyiPJGA9pe1KQLKBqkBqmmt+DDj4EoegU
DBEII6FhZLlmGq6uk+wN5YMm+XNnSRhZtMZH7Ccgw5Xwub6b1mySb+jE0z001CXiCRgVw2uXUkTn
rg/lBAa2te99FvUFTGYevUKigwpDZchdNc3uhuecS76gAp6rIkID0W6LwK5TKU813xKcvvoIzm24
mZnK83hkOvgabbrtIPxthyVpzlWb1vOmBS6Iv7nlm697rf3T/ZQxXlR8Gfdw7hlwNU/qlyV3ntON
3+u5O+h6wSHA4PZF5MER2DQ5QKL+7+bruPsRh1OCJRyp/DWRIBj6t2axfQB70sJuNswoxSLADdLQ
ADZz9yhkXHtRTh5aGcOQ4IA7sTwG7EDSaaSQ+1W3hgJnjhjKjQCLGg+vS93QmDv9RSPeT6nemQ1l
rQvvhjQt5840kUVJ/A93pKAj8b3CP6kg7L3n/bxgxuiq0tWAJB45bXic15HH9M0/79WWTwLv74zv
oZbCdGDHYd1+qfdiKzhTn07XVxs1/3WseDq9F6d9zx2hPjamF1hAvqWEEuabrEfVy8go0OEA65pw
lEfr7Ly7t+FtDWpT4Yo8oCphXspMzLC/TydaYIy9Qjg13BiQpkidIiiOjOOGpL5EKYknIae9IsKH
GP10jvZ2wYfLH1aGtJcReZWFFaEnq9X1i/MA6E3dRDS7fGPzKvvX5XARqliQySoBxd0zKswz+gwY
HqemYkoC6V3KiDiz0HxW6XINaDBx5A9A8AP7wcEeTjWE4nnJd0a8kRXbMPCQ17BM1CgI5kVl55AV
kWil2iR2J1QRl5XDpx8X5N8CvbaZnlHsfIYgji1G5MGClK7+6+XT/Z9G5wcwIIbAUfMHoFY9T5QM
rS000OfLnqVzN9OB9ob28OvcJBWdxz6fli6FjFvTu8TmlRgk5KqO7+WvyX+nXa4WtnX8LB42+NFJ
owbOO4ucbPPzvk7oNBlAJIJbIiHgZ6gHwv4OD62eooVgk4l1tWoVxrlprlHhZqeSSGzOq2XNws5D
PhedftN2iJtLiLPawr79qUthQ+9zmpX59OyegvPFSakljAF4UEO/2Gfprw9Mk2Ss0jho0bN5w6zx
YoFDJuApTE3/Bpw+dzwJtPE8p/p+GbJipoGJ3MhqlkHvUbaxuKhactPy8khBgfKbsDdr/iU9eFyc
yqncV+irXbBsP04UkCHp68Oeurv0Strv39LEPMkY6A5668zlqe/QwcxfYURgqIdv9R9jqwU0j6ze
GaruHJL5fGeWtslOoNrBFAL9BqutVLdR8q5TsINQG7YVd/p36X9Wmoomze3SsQosvduVYAjAqm4v
25WDDOCoBjlvGmXaCH+lYUM49yM0IXVVFvI9hhd0Cfuw8FuaGLgkhCmu2AA5JnJEUrsI0FZP9Vts
isQAmcb01bBMQVrfnqo2wwBSuaMRWLTDK74jCYwgPlGgP5OyMbic4Zq/k8zkmJuefxQsYQNhk6oj
8t0dkd2pPDmWV9Py/SmeNsAqMS49v/3qVQRRNTvFUsDx4Mhe6992LVcceFBhuFjD3te47G7mTBe3
NWwqO0SSMUjTTfO5erZPZmZDO3N2dNEMN84AiL/BCPFtK6+xSEW5q/YewSesbTponPPMDNJN4Hsz
h6xkQBIpNC/jIWesCsRkpd/AoxiolEClYz9zviDFInNO214Z6ZuvPCYwvgnd46yan0SokxYvv6YA
7tBmPl6plWBTtSzZ/KEYD6XHH5lHYo+MeaR8SNtwEnwmXaS83oaoF4BySniHPbSg66RPHpNWMrkR
JOf4iJtKhxkuovHnC2pZyaZjfEUpNPvhNKJ1K02/VI+XIkgA2w8j9ivYqaFubbZZeQtQoBFQp5wD
cg3fLEs858KyKX1iTZKupVWtKpqSlCJtl2LoQKPxutq0rVPRXk7IAosL9G1EMi9emjbYrqk0mI+L
gT89XknNZg4Ho/AFEut0bskPk6/NX+lT6/BNMjiZmbZLjn5BwJEhvnJN/aMz4z6R+r3N+ZqQlqSc
6iSGyslxEB7lUjbEB9OfHgNc2Z2XE7k1n3W9tCMH0SincDJDyrClJmo0Hn1miYn0yD2lYFy7NPci
In7wLJWsrTbd9dgdofz41ZjXXj5wIBtCrOOZZz/FKHfGKp9MCcI0ASqOv2m/cM6NDxLPmoRCc0sj
2b8f41cjayDOffwmBQZgSpcO/E8xGIIjzKwngj6JUGEclt1VjgvtKLQ9sZPpvyhczL803S2bMmRL
rZofFxjRfh8s1Iy/fnFVKz6ILLabsYQ/sq3SEWErZu0/1QlZZ3TelLzlX0lXshqK5+s2XB2Ca3Z4
JFKdmNBI9KODBZVGAOOxNorRYfEQXsxQxgRxIj4wNM4J/CBvmO0usf9RFAuSjK+ZwYwUUj7dJqZK
4Plh8xFAbuwy3rqPttiRaCyXXFQV27nw6J/TcnCB+zYaZNKdo1DBeCCl/+MZJ4/CpPbfjcI0avZn
KVBoqQ2jAMdIboS4ZasIRjrUcuA0Fya3zLhj/+tqQVYBEOBUh/nZsYdzazFjaP0Oh2aXrIxxuPP4
DEcu/y1mKfMm15nCHzSS6sNoKbn9X6FKZs21h8EAJB75j9EeOoEz5jfMA5uTFxck6EYZjjDuYbva
zcm5bz6mbSp0rUPM/0f55Kc/qRiVkj20KU8zjF8D+5psMhB7o36rd/yS1anLcXSs4iIXf8TKDAVK
/uumBGoCDZbcF/qybYqn2b1OKBljtiYBEom8xeaoSS/X8MtwAT8XWbSuYI4eWhCTa0JUfKubRVst
sDM6rs5ZbpoNDQvtUUWcjLp3Nvw7TC4dJjP4ofMHjrOLxbjMao+OododX/+YvXcxJTUiCk+3dznX
oBa0ww1KO6wfqilIY/0PZQwb97pVivFo7zhcVreDm9Ry21Un2QDL4jRKmcnOkIfkjrYj9eMP9quA
5Xl1arb24NnesIxmEtfUPvPHaFdueHXonLLLpQjR/MtqA0dAcmuz2k1q80BJLwsm97DK7K0Q1yhL
bt3gowH52iz7bYF8M/bIuzQ1nQxLX3O8GmH4ZkM+GHdo28iV728oqiQWJPaRYQF3wY+V2uDCjtK9
D0rPQWU9CkGoCF23P2H0ZCNSZVKU5M0nKAjOjEBjHFYNAYYrk/EDJedxIKTbZaAMhnHxS8yCngVr
Mw+3qpuyVhyN05iGVakGMCQdtxDWhQPCTjL3cllScpeGhVHZfQJM/sKFjnB5xg7RaALGPEz+I+qk
2eB2UAWJ7YNZ4BJAwjkTAp4QuTjSWzXS+VIgkbgaJswT1GMTQAd3llx5NzDmEr0SWCKX2iHnQ0Bj
paSY1JeXWuFxUjlw/4ZRFQGKXN+Dgja8GU9QJuN7izDTzCHFwdvqk/i8aqIv7rGWgCk767h9WhAY
VHuCYNpC4cqodOIZxOV0M1o4INT9Ald9LE7ToZqMto9aAsx730Grn26GLcP7C5uFsHIdfxkWh8XM
EXFQ/VqzTo6pi31Mv0H2BrLjwYRBoORWu/B/Lq8LA1YIDEoGzcyt0udgEbTITBvMEoCY4W8bmj7i
Qug/vBolgjpgi/uCz94ckfcRxf0zJ9njOGqzK36xx10XvaLo3mUkiw8yyAcMeJ7dKbP8hzJpDESk
nwd/NN839CEEd/fegBvjPfctZHFsbiUu6WABKxnlYqDfckjx+qaN3QKYcM3QQh0+SC9TS20kibQf
77hffJ8dkzypVBXn0JVbyzj59n8NmPIIrv/LRtr80NkooQY/z/WyJgUGAaWiqKppWrfGLGBPNCzI
jvwdL1jwcAoprUrLzPrlDFpoNS2QHzo3wcOqYg8p6WoSja4Rd7SOvDhAI5h9WvlXWAxrhmlIxT7G
A+RwdGST19fAg5SrmMYKXNWUhYqelogxp/W5ViR5SB0/8i0xEG4BGvd/51Bu5GRLPMZWqN1phfj8
+ywUKOHOD1HGGsvXjxVV5QhrlHX5WF0z18sDXjd1Z9Z5PQdsXAACDkibBUbrpH1N9aUNOBi6ifAy
Nl8cmHgBEZs+Ooo+SNVaN1eI9D5/8J2p+z2ujkPiJgvk5BD9dKyiAN2n6nL8ESZ0SE2MKJ8UUM8Q
wZ2Ll8H7QWFkdht9pC3BFC3a/0CWJmOL+iB1PfsHQUQC2XikWKWCywJ64Gyfoli4EKfabJ0dHR3Y
AAibefOShzdoE7mKFXnJzrA+mx8HC788xtkGGFtxOJDfmTcbmYua2V7fShEGMZPU2GgZq6c+h7jX
J7VcXabi2iBJQg5tTQtf+zRTU5owLU2Q59n+6pdtRvXrUgLGPHgdW4fa5UFA4lhRbPZQRb0IL0ep
i4Fo1rL9GnIX6EN4jE9veFHpxFNJX+cRqxE/6QGrTZyfQJ+XcLBkgEFFtm+FbxxgIbY/gWj+kPbZ
0QIsCOwKS32CXLMQjWiw7mb0dEyiXBGCfEW9Fo8z8iD2JCqVEYEtjjVqflpgsqbR/rhI2qKVOxp1
m4TqMzNAMbEIWo7BPsgTqt7dbUktQNa1nxglePD8kuEOZ4xfSZbZKHITTr3q49tkFtSfLVglgvoz
lTUgYXefRbo8q2ROCfsNfIagak83KB1hN/+OB36nti4wr4bBkzDM/GyKl+VQDfu6MBPi1zBplP38
wGhSpmjggWNrHO41poEnkpixpqOBVj9co+qB8jznMnQH2sWE7Ko3NtsPr1KxR82HWrq3RcC/uPoh
EEt1sdQM/yAeZLwNF1Hmb8J4DA4XWxNDjpLqgE6YNGmZoIhI4mUuTHwQEgG8sKml1I1lNh+GPnb3
Aur/F2vXWFwf9ucsWCtn2oLjJGZto7WPIhEvPR9EQNOqdULcSE9XgfYPhd+i440DxmiYgDkBrm5X
N4sdBqOckvvvUAMs6yRa1psYjBdytmtVAPMbBrkmCIvyy6yazRvA/XAzmm15rhbOjRNZ1iAwvw3F
ipyog1YqLIeiXGgBGUNZIYglMP90PMUYy+BLSsLN7lAhu/qWWndbMn9xeazaV8esYhoH9N/Ec1Ij
gI0TsZ9vbBBBsAu9eEGAgZmcFoyZ4Fuq0U9idlW5ICnAAleLm9etjBK6dl3XjHhTu1elOmhl9ViB
BykRNZMUsOOW4KmUyntkB1fACMsYMQfWyho/0smKPfuLldU7JNyNE24/gCQhaQc5lRjQnu0FLtVy
J2hjOKGCbHqUoGBTt2eD4kK5EEHKXv+YBOAG7vOd2v7zXxfaeRcI7A0vANbFsvv8rumnhusQjFaB
w2p9ElTkkcyj0/lnNPMrcXfUhc1dfdrc1iNMVkRfHAkx6hxBjCQQZDeINj/kWQtt5wWeB1mWZhuB
3JglcogmfyP0F0102KeZvsUbW85eQ03QJFp6RXuEfNNBWzjxRbOpKuNNviweTJvtmicw/7G2hb1G
kWIyA71TGQVryJlonLWYsRTgTOIHje72cewo2SSXGxZ/UiF2PxnoboRjVFM3b4CF5z2+vLeNCfRh
6V8nGlJelQzcy/Kx0qCItb6tuhLdVG7aDqg/jRo+hr8lBzhFUPFuBzRUQw4zE90NdcE10m/CUXvJ
SG3J94rQNTwz10nICMp5czulaBGXxybZgLZ3xGOOzVdzEidD6BBhy2/4erGO0kdhbqlOTsqXEa8y
7DUg7sMZmuiLZVc30hifnHWWHsGvEArZgluoHjL+ccdzbknQ6MEbq+3b1V5pzcU5tdHjVbkvruYY
bNzZI6ghZhJNO/SoYHaz0xFtSjZf5PwPzorwxLdlACL1jsO1jcSv0LijjwojGYTE/Ihq/PlYMSQY
o7oqmbXM3hldXeKtmC1obl2cIpf190bb4rAfpAEwzOSRpgsejc9EmAQzU/dO+TYGRY2DKCdVOzhH
27VpugVtjwm71WEkPEnWcHu6vRk9oQ06xsNxuu+hEiVtDAaDFgL1VRFjmofxb9875eXuWK9S2M4w
Lw0YSmTVXrPYCaNr5joUxbJ3sLz5F7gux33V9j8R7UYR/ioOrf1ET7eBH7E/X7tiUZ9iBudUWDrM
BPuOBZKsTmFWnxHN0RuYtG3jLcSSvK7xLIhqGGpMHsMoP13pRWDYPuRJl3BJDTKLVhW6gt0Ikfco
Ey70Ga/FjjBsIWSxhRb3MpcAxvDwPHJdUH5WphN4hfw3esXpJCNAVdx/+o0uqRlJGRCHKb/FO+YO
9rk+389ZHsHUGGmYqREPr76SbFePL3n2LVPnPXaeb94ZA+UxuhyCO7r/BWYbYolLMfwKIA6NPIKw
lKm6PYLtEJceB967o6zM3oQsrd1WiXEIDYZ7pbBPbjiKv8/XuNOpA4kcdQxa0+YiwRyMu+JtMGqE
CXyOoHGTXHbhbNjMtB0CTiRzlBw2/+5+ia3LVLyYFGyqwbyKDmhm6+GC8SKZRu0PNCqL9CAz9Pz+
c086nbnTcAa9RQIhXB6zuxy3yetXdJKgNEr5jJmZhtCEfqqWLcuBkZuj93RcUSTGEfesdrq6gcAg
rOKEIcN+s9mhlOMmHbHSPvV9m3/ZdjU+G6lyc4hS7wLj1fQs7Y5V/qejy7pBiW6QY+7hIXQfTMj3
wnyDegqLLZtpvzHPG6sSjggfQx5BtrxIWipQLHhR0MsPpCn5Zoubp1fvRJVBlG+QDG5KIkhUwIjY
6ViocjfPWFXjkJKrQl2Rih18ZujN7sOQ7mdbAPw4JLsvsZuN6m2udtQ2+iV3nJX4+y0GBRimTc9D
zSD2JaqeMSsZAhmVIWXHviAm/8LPCJnObcACYkSasMZXNrrU5hZMfn8A+IzPmlmN9TEUBu30cmBw
cUTVLtlgKYsOB3uHtkT7EhVpJWnxFrm3oMEU1Id9jujb+xwPjVvregfbL2LeMIdrYpBG74Y7jjS6
lCLmPOlyIshE5vV3N1RFoxPgRq3Z5btNGIV85grgxVvplj6zabaZp6rlr49FVbN5q2RIEmtbMmoE
MTa7y23pbQTD21NCqDhS16N/dpQdvb1tpsxzaz8Y4eza0eyFT7L4vuC2kkI/dedShSPhE8eR78Db
P8L0FeMep/nS7ULXUiPAzdHWFgj5zp941UqpcmJb6WsOqhk2O6nnswsZOGvb3eLe5lWyLP0G9oDb
hlGe8wMGOt7ZK03Xf6gq0GbGOCmAuvHxOvSEa+0L9s+ranAo7ZRAqsrdfGmglYVTqW/OauhKvOWH
d9syR29qTDjyUFn/St8Xr/8ZF8fLPahWn884EPmdO5RIBdHdGZTSV1asU+MBbLCVgpQGpcY1eAZF
HU+h6xGa39j0q5M52hf5NKggiqRTJw3HZziy8FdX/DW+Q9YvMLE1AygUTt3qw3/xkLfqEOwN+Vbq
VmaHQ6rcYg3HWReYndkN1RXCTvS/+SIh7f4BpmuwtoSS/tN0nZx05lZ+N4Dj+OREUiRiiOast128
gkS2UZy9ytNdCyqnxDK0iRirY/u9YpesMZY+Q6YidG9jl780XMgwLdNdQQNjhh1GFgMGuSkZ1Dnw
v/tfAGcoszv8vVU6aTBKARv+vkJfCD0a3h7AHAF4vePUuKmstFI+D9HpmRjWwcb2a46l1kog9KGr
5Oe3nIDZOouaScJ1PovRy0+fGGXO74kONWuDpxp7Q2a5kKMMwysDlc6drqNeRaUQu0u1XoYlO5sj
Ncf5/njQhlDgX2Uid1iwgBmVk++YtYg6nqhLzMt16h6KVbwFNXKL66z5v7s6QQtzEgG7ywxPkRtL
GhOIxNx5QTaUMaVyE9DkNQOe8Wn0Nv4iGhkJ1qjmDhwmRK3j4J+JKmYqG6L4vIGbFQzVCkGIJhRH
o60ThFy3GN/aKhGPSkV/FzZK35gJ1+Aok3CB4WE20gs11on0534WzBFdu8QOu+i3sTYvlpX2lZhs
b3PeFhn4dCl1MiB8JR+x3QUuC2R+Cz+6bvNWBiSQ6El0uXzntURxH8yUM/UZMXvS84HBLUvCZymt
1mnaOdZM+Zlf9sSSkw5a/PE5sImFsPxhYE5tg0Q48mH2tUwSAKPISXn93hdcLCOrfO/fnBEyM/+j
nHuplvUzrlIwUy6y81hi95slDB1d3ZqXvzJuE7ui80rfZM/pqczbwOcU98S1lus+uRJX2tNG2KAe
SCMXfn6Nl4C1Fq+ZIj17t/T2BQU1CBUafxJGVzpaeUiczdc+hRz5//04pZpC7nl1nv90HXzAmVNh
Ek2YslA3mtEL5ier71xSL5InopXmxkOk3RDLVZBf9Dvtg7SrDq/7KBXFNmcfZORk1H4MnA4RpL6W
ywjdUMNtx+TiiB8y6shDSS5Aiqnl4JD7oi0Q5kot0VuJkMQ7XhAoGo3934b7bWQG4I+UbIYR6sC/
LeM90lGzKEWie7cB8Q3IISocubpswcRunyQgB1gMSMhZgdwPe/nzfYxeFO+0ADbUXQk/Xd39mCaG
TMCvfFCD3obw2Alnj1FZF4Jb0WPhReiqCeHg8jEiCzZnJEF5N4jG86VzKH6vT+VBFYtNhI0tGk24
1ZTCbTEXtX30E5R8pB62a6XXMvPreUBEFu5czbM8bzWJYJJe4c+e7laE8kZsOX6xWB6BMR3lARLw
1qDoEknuKA+QFNrg9A+t9SMnyJipH9iURxrYwluRWI8jtxS4gco6C4f/8nEeIXZX0WXLXGm6uUFa
beIJzbUCE5DWOQFM+nv1Bmg1KS5HQXXE7lWbS1Q3D4gf0BleBz8YKuay5ZXStozWvaP9aMOWLhZh
Md/bsDfvzhX214Sx4S/1PdjLtbP5n03DEd4EqZ32gx87vv3gNaumaeb1p8/J2te9fyxOd1W6G6QQ
msWPRYCPutuNGbX6XgCt9jb3Eg0uB6bw9JWTPXPmY2FCZfj31PtMzJbGChsXgJjHAv7Yp8JsK4Mw
+Aip9ecTBnF6S/Ezq6NwSm5IQYjYhnq335/lOCa84pAb1xBFtobZDhmtzyq77v92/zLttnyZKcZq
+G5jrA96s0VgAj5KB+DK6n1GO7/pc7ggWKjDcYuMP3c8M4xakZ9Sa/6+Mpv5cJVFR331EclY/AdC
USTv9sOzhAnJXvgtgdtUPQutSDLhLLGijjjhuTSZG79MLS9xAaguPZLZSfnxGjS0TNHLrqK/CTiW
SDyLlAqAvJZgKp8grwUtNM/2w/v2MZSN/yFZJmFHMs0QJ3/SL6ar5SVPQA6pDwr++Uejd3KRBJa+
qrJTc1PWR/f8EgMz8u4eUDqlkYRM9G9O4B9M/Q39mY+LwNloAoqJbK8fFBOgtGzYvuJlW6SFWKpM
Qf5Ma3iEGlVpRwSTF6uzZNIU0Q/LkGrCyRbeDNswzE0ilLvz2ghpcMwVQ5B7OcaDcxtfq1Fn4Nz3
h4yVMtXUJg1SBznK+7d+/7+XMCj/qZGer1SiVo2qJ0yQCjibbSHI9jKV2ERLcVU4SJJAwsVuDx63
L7vdhVcKDdKtNqTc8ebgzyYJkr9/WML4r0GKoClxtTN0onLifShZFP+Qp1833wL7/MPRcU4TYTn6
TaNgwCmEmihidJ499+ddmrsu3OK6GL6wRRV1kIHSWCJ7MZABZ8+joaxxfrflQwOuLVBtZnjceuWZ
jXppAKdXY6HhHw8pfmXXU48Vq9+3jvYTn8fOyK3j7pFrAWkWgngmIYDoGZphswdzWVgRMytIz5Gk
J07x1ESPfxFay1eOF0/01Rlap/EOXt0VtUBQoGv53FY67u1HYFgfmkNJPhdYM+s2tlL1SwDBWakg
AC7AMQSpJt3db+7zXagjFpbWE9+WpgV1VSwGA1THgq3rzKF2fCezZDdusiyQvXmqGnDb5umdOJv5
aVccMp1n45Vza+IUZ2EVlubs8ezIOO36LWWRkDV7Wa+bcXw9sqzUi8oPTYDi/Eh1NEWvHhC9gCuO
Ntuuy0z8d93pLqwluI/yNYsap1TidyZEZO6r6yTKWTFYUfrMTsFRZUqwWJUgiMQob3qSiofjVIZe
0HuLtshkDmmZ4i8HqFxBaAa7Waf3xsGskex6MDqYOstLLyL/nJ1Q3jk/MExhQYLt4oz9A92uI9tN
zal0ONIQg9+xVGrUBjQUjUiKNZxOzOj0OA6OFc32YC5sRCwX5sRryLcWPl79Ltwk3WEJUi9dBUbP
X+m24aRNY+gsk18JuNupeP4m30nKFJqJwME8zkAGgOFXS4L3gypgLA+qX7VVxH+iQUHPXVYC7Weg
/hXLVTVMMc7WCBSpkIrg3/OXaJ6fs93Xsk3dIDAiv5P0E/TbhuNFOYlNFNKMMxj8KuSLGIM8cRmN
jxaox0UVroD5ikYGUFNvRZXs2aqFgdPAPFtyqhkP8u00s6FdT4vPCaJ+MRVBExEFWH9x9He9th3v
tXsHHk2mmoPC97zQextSurhgP+8NghjSIVN+uvuOKXroVIgNehy87CXZZs6aH3G/1x52ui4YS44j
D31Fw6Vf37YM0pi8tREZ9VHItphL63Rl0uJpwSYcV2u5U5RUuIZ4Ua/bRWbVpCrI7mDAzxTyK7JM
hVX8k8U21bsx60J1CIzLRvrQRztdsR9oAVObznWTSHGpD7BwZd+TXzPtMJmqYBUvPiLbFwVhEN3h
4j9qDTUWOd3Z4uRunXc7G7IY3/WsjuyuevPXvhhU6TFQNX8J03JGSTFdZyP9jI9X/EHKJtGr2WlZ
0hMujPpForNPQGrkc9IqpS5SMpEV+vlSHSNiRVqZpbpCa7zaffNoDwry7mZCnJSp678Be9y0gjKv
vp9LRHc5Prwsd57eOIPubkPAzx3ku38ko4IUtvNxt/W3eNS3+s8Y9E6WXQl4Aa+25kWDb8n4opih
Znn22GxtE1v6OTS2GNp/+DD+ghefYA6ynyn4bxtnKcXSBDZY0vBolsqTg4unt9OzgdF0pgKrOvEt
Gw2hmbO9L+j9UTjv9tsy5my4YNohlKxI6DcfjgsHnC2W/yJGZXo1J35oSX8Ino7UF7Vnh3KUyD2e
d5K/fHb1oynyM2AgWmHA8srXj6vNEiXRSr+K7ZRGNDU3Llzpx/20mOoOfP6LSc7KfUzceV9a58IT
VoO24IVqko7JsTQAa4Nghi2Y/gGtkPeiwKIYkN8xaqZaHexnqmLUQ0CG0YeQ2ZBpK1j86oACzbLS
03nw1L7BFPF5CLfSdsKicIOJWyRfCCG8HsjXP+KcVFmO2DuFp41NK7mk0/CkLHzu0XeX3Ro0es/w
npN5bpEoZhc7l8fg4mK2JklHvgg52a4pRPpj5stGtjJM0CCFXZwjmSDQKgNVHrNGrq8putMfoh2f
RC0Q4dZ660JTydYppmUbp8p6t5X/I2oi4qj+rZpKrPF47Vd+A+Zq5xVormqhC6juCR5qdzydDqdC
Ch92LukzZkJR//DuQ7+eVJHiSmyXFVDZFQRctGVZRr+ia1NvohEwOWIDmuiGnLM9QjkR2wMz8br7
1EpMTC1Q2xzCIcEpnttngGVz/XuVxQBBPhbGJuTEwxR5zZn45UcoIGTZxB84bmEoXpHUJ6lqhXYO
eWEOnenopqiH5Ap1BuG5gvztVEm9jbb/Z0pD1c5ooLKle4jcF3Z/xinDDpXtoC/+iLKKFx95FyWP
YmUA3tzVaswd2V36zu0fCfWRgNRBlgy+vH1mYHn1xY0fjpRL58mQjT1d8wYX59epXI3fKuS3GyZN
nwZXg4VFq16PzlqRocil6yi9HmKe/KFd5noleUq/737tccLICwsgBKJuC6rjNFd+6wPH3Emn3vXS
W+o/93+zE82PPcJPUu3v2QDaVczIpj2mRwCQMR5f7PSNuXlsNfQ0krpHZqxoXnCP+YSfihaCowv2
VlHKlBrkahV7vqv1bQ/kwolyJGZ9ymm399Sw7QLlyRai+Z/6uWwGiqm10MUSmKj7VWHiSARm5kTb
xaRMOsDfrK7Q4Ozm4hwClo4Wj4tFWQ9H7NYlTLIPiRwrkPEBfARphU0vbjo5CiHWGGLmY5xyTaQw
5sudgDMjJ4USMEa2tHRs2OgfH+kSEQPeGBl/Ln2VTCrczBDbaHrGWYwu+lFjT7L8E/ZG5ROxScnx
TKa0RgI4sDLvR9mgyqe0XY20MqgWAoelul+fAcb3mdmkAGyBvYe8WAQvyQu2RofUTQSAP0LvVahr
7v4roC+wXSVbLp0S/LFEHoHHCbGlZ1nai/fc/AUCsilOSMzjNbMFaS3Gr0fIXBmIXM6cxHpvmJdZ
b/YYXUMRd96fyP8ZJ7sjfTvf061SG1zvdfNG0xjWBCiX9J9cOTIIEsxzbxE3Nny/B5bBx6VCjvEg
OoBaQgEZmxRq5Qiz3OFzQHdoxbpfEWWUO14ieDCJ6lHQ8baSivW48AP1wdFyDMgGPjD02WpRiOx3
JzvB4jECynhwadXhLbWTWeQuZ5bxk29pu1P5c3MsEXTYfoNxQmYNv/SLln+6JxqVtkKLabDtgUdQ
5Edd//qKrXbCVq/ioZP+7vfGU9kAKiqfRsa1MMSMjBLLQQ73yUc1J6dG0tkrSA996EL/INKLrAgP
5ZqD5TzXYCj/g29yjtqSMTj+TvcCwuk/YG6ZbJYirlXLJs3PILU1LAL34fSqtQCI8ZMHtGVBpKj5
5HXvv7q2RYI/XsED1IZ9V6gnrcnreSbRpROIlGlug75WYD4iRG+fB2ocYE9mCLVxbDer926doNbn
pr1IbnycUarH9vj5lUH7uZGQ+9cCRJh8f5GG4pFpN1ahPp37oonZEGfL/rRtT+4Bhk1X3La/3D7H
rMn5L2/ymtWfkB87IvqTeSErVAOOX8yAl/3vpQZmVIhgTTV09v/NXo7WahdWEfbIi4+LcxqiIZiS
Oozc3bdnnEXgt2NrElG0/VIkGAI7kNa2Tf2KnSgjtXxpNBY7zLB7HW0Tq2cTKMocLfQRX9aMLv4Z
XLVH9ArsQnswKbmUKkGJGhXLGtKYgUSC4XuiTCia9/IOTFq3bNXEftwBg5vi8ayCkF5bQi2POFu9
ZviBiIgEZI34sDAAGTq19UOIp7oBHk/AQhAmcDJ4XlHrb6f7IOOO7c+jJ3FVGdswO+1i+8hUT0MT
Duo+EZJ1dFgelsSPo+Mkifx+w+Cm8+y902LEHjuIwPtyFXCSCuFyVZQvr6hJvg4gZfJ/eAtbJbnZ
6zOIsR+bunKFpo1BbU/8poX2i8Z/hXbD/txYO6cKjBb9ywrQ47Pv2h2JG39OeWXpA8A4zCYtvnw2
S1NxoZMcwGTAvx8boUqDFyV4LDorp1bU+/uPNvr7vcEGz+eqsY7a07Fyzid3BUwgPsnIgaNnreTO
HGbF10rhnbJST+M3foubKIXbphHUN/cTLu853yEPAQ7shMMRpPqQXIuUIYDQZVJiqTj89u6h0D0p
yQK7FmMqqQ/NiiR06s0vK0t2TSml4gkHeaxIB0S3zhZYLE/AkHMxmXqE+NSOO5BGx620gPmti2Kf
fPK6+YmgJV4adt0GqmyqJV8jv3O3taaQNIVaT7GJlUyaqgOSNKMBZWEolkBir0WSUeiAzDJGd+0y
iJO2e73hUzSbaIMCYpx+pR7uizVQzbVyntM6kw60+C48YGbMFdLfsq0cOm78f74Y02XHnYzFRc4P
mY7QsAVu3coymYRGM1tv4YVm86hzhL97DaEGDPrb32qhIMXMU+UB3MHXivYeK1zw4R7Nj8VL/wtu
nrENc5qpAe9VUwPKE8q/jURP2yZ1C9YjlrmCGAeC/rmLcH4FfKJquRYxKy+NUWgLFZBwn/YL7uXH
7/KEgHoRdey4sqIGd7Bj2JtXLiFq/Hs783rMA2mW1ZLkzpM8NeprYRrzVnA+55AalPvPUg4b6pfw
Txs0HkUivXSBJB+owiukRsf49GQDVUxnFUF0zeQi1YmYef/6ULWDgraCQedSei3CctP8h5TMNEjG
69UIJ3sk8LUuMBwDL56XUXrz71Qayxv4PfsExpFKXdapRftTYHcWG2bbzOtc5qkipcu6ZYNqdSjU
yt6uS/ho8cAHOGlkO8x6rEvd/JawOrvGLeRXb/GPhLWaeYHMsfW1dkX7Vz3AvIf/DfZYdLxnVdd7
whgNdOahPVEvOFOgDpScywvF4+f90LebpVZ6a0u9mFg1snrLi98V46Q1dS5MxsfuQU6tFwkVyArC
rm/obl5MuchY7lR5xj/67uUFYhEg3FrRlrH3l2oAQ1msQw+hCFfv68cix+EM9xMSlXoC/FnGHHkE
DftH+N4WjMgOt4HDyB+KtotN5xA3vpcmrUUYw0WI+lvLrGWKjGGHDB1AVywy8JhGqX45Nov+ExcO
XxS8mxVaxS453a6XhTgh2PD2g4KzW0gHOjOyTcdhcoUW8Xj2UIP04jFz+Eq6Bs8I0fvaHjYnl24/
KaYBgYbiq24d+VmCSFbleOFXKIaRvICegBlCZ3Yg8ROgY0MzeDO59b0A2V/QWlQSeS7OCEYZcHIQ
cFKWK26o3bS7Eo2yYWNErOrrw3WRsQkY1VR3xhm0mYKV69ENwlO/BNGf2gpVdjMiV3wXiok7Idy9
dQ0nXDqN3lt9C3532m6XhXSpbfT56fcnYIazD2NXNZ68ffgq8yE21sMSNB7Lo52qBiN48GQiHWhN
1Jxw1evuMFK/XC5fGdeNGg0XVUl68M2ipow70crrY6Zju69UP4/VAi/gmou5mmFsSKwhryfXd1FX
ulGDJCMoKS6mcthLkkZAekj3Xjewy7q01u1vSFohxsVOHtjAQgndecYbOJkr/XBbQiVMCV+d7CdH
NDYbtr4Z3l2KpviwlfU9vRpaz6ceaH/hpnvH6ule7EKhSWTkhBi3sx7j41w70vOA+ImPfyiu48/L
yGb+QpzUCJZtWpulg2PhbLELUiPaWwqH4VO8lIPUXgG+KyK3nTvjiexlfv1sTKNPTMzl5BSzQuDB
7covQKjALN5cytRSuhprhbZWAsy9tPAdob6dY8ERkhRBaTVzHDJog3AtmtumVT6zwA/FS12BR5F9
U8wRKdKeYilelBsRFtAriM1kzI/SU17a1gO6qUxl3Oy0LRoTk9SEX51Dj22l9ccg0gfvYRe2WOgM
ECk0aMk9TR0RULKgpkU3dmb8GzuM+jFadz8kzo9pkokNYDGz/ydxo8rlYqm20O/6gzxaxzcpIA+V
mzLucyw7ExZX92AJHBSOLSYyd1RgUU0PD/lP9TgOYzwp0anRQt/PRZ2bnNuHCl+KolyHlhbtWspK
CwK7oVZq2yG9ZfBWQdscwYqmTiMI/lo9LVRh4Sad+IizRS/Oai+zVNA8WvuFpxftldJf0D9LERI0
Q/IzOFNjdW/g97n8xp8jlzNJOsZ85dP5KYcJRLHpRmE48+T/aWagj0FWos6jz7mJEczhTV82WWEu
75E49vw9XF5uzp/PNtv0fG5L4Mlr4erHefHd/HFmKIFqL9Vn9mwZ/iHJDIQBmQC+7tg7BEXfnFLw
hGn0rmeBJ9X9WBA2n+z5IEbz+SB9iKBuAXt6EHugQ83QenIo1XhCotdTydApggejO3IjFip7yW6j
x2/B+j1JfnPJgfE1pCPXNbCWcvtZMh7b2cM/tm+DvQO/viES003A626oXNHVqmMpjKrcwMQe2OPx
hd/sToOtAD0xjxcpwPf8V3NkWHun/BD0KY/UZS4vpycQnLDzrTXlk6h99tjRg+BKW/tV2uxoEPjn
6VFrjkHa0fokId8kjLmB6DGz6N8ZSKmzT+Yr5B68cOMj/1409vOfjwFNZHK+7yawEAMBO6YOZpaP
CmYcMvkL9Fai9J0+ctGfrvVXa0PBrTFU7TmMRIM7/xpkruv3BiPLC5u8dxZhMXZKnPIrPc6egTvx
Ky1QzQh32Xq3O6xwObZOMAqwyQeFXVO2xlvmHvWsehelri10QV8PLvC9p/W3C2toqseN0IjmD/To
wHu24fuKo0mKgylPD/TDQawmkT2QAILeasBN/ctOujSGt6u2Gfr9dVqtdTNt4mQwdbTtNTXxOM4f
okVMBlUMD26PCioM4RS21wJcYHeC4ziz2mkNZ4IMYiZzFx9QtYL2j1iJus/iMeYF5IU5+XiPK4k5
X5z09s6ZYYMQ6UBkXyMkm5cNVuNtOrR9gkQoiEsQAdGuiToRTXw+lw/H+/CKePOkybKocZreHpGI
jz0Jfo4KusrnL3uX5gsl+2L8wlVYj9XQG4xzjuUM1fG0OJ7mqjZy8vKofUi1HpiQr9bKlckj+jfR
m3IYKX0vVTksvuDopDjG3M2/AZnSBDT8wZH+z6cms1AuLxKCAJxemz6jOHvhgZxyrnBIinJLhkrA
H6GphuW/YjY2rsGXvcAQpDwcdvuYjjv3AwkLTYft1zI3Gh0jot4pJp7EBGwq9ERnO7AaJZa/h+7f
R+kVrJKrUIvQwCKjDImIvuIwJdqgXADgRlv//NCb8uDN6MELAysfGYqAsKbFLwx+F8c6Gemle8vE
oU0OzVzbLuLcmyUN8frzkYRh7vd72zkBVvCgzaeVL1xGiP7zSUNuaRMoK1l4lm6bMz1MJ/z0flBW
lcpA6qrDPMwPeUKYGRy7y+VYPkxQ5NwqvuluH6gOSiOvcSqE2ZOlMvaynxq1tndkMxNCLQLYgKmE
1uTyTAHSSAKGjFklJQnaLHNAko/Gzf5oajFtjSq2C1y8E73CGNRn60TKL7pz/3GBaitMnZ7/8IwA
4faFvMaSdLFv82Gv6yRk4+sWAqAaFeHttKdpmRARDOtEsxWSKs7NPxyTddpWv1kfwGSSMKEawQ6U
wExIpFxObTTybCpU9LmRKK6q5WJBG+8+DiN/Lw+drEuSygEHlVdVf3mEe/+rTC4cf89NJtaHx3xD
V9+tI4YMIAVdU2cvqsk7eoeYv6LJElwLUsBhU0cKmYaSHidkx3vj8ZNMg714uRd7TATnJNrhjzMT
EklreFRWtgWshn9PUktw6BHfZ/DCIcntBHHG+HnpWibJMVK71glbLon6CmUiGr2JZfukjvAXqvun
GkC4s5uvgvcRETA0tBq33OXpdyYkp5L5ASW16dAkNLEOLnfixPCKKf9SbxdjB8o+Fhga4UkHomCC
Fe+NE8A/k0jPAXocKZj0XOAL9WjgzxgElxznnq5ChNrw9zyRrhfXz9IlHjt4hxGJmA/Jni2yJYNd
wldD123oZzwkcGX2Lq+EkYxtQg7XlUv09lxbNgQXIG2rtEXOK3PAS1YV7g/WZ68SM8zXntbutFeB
0WuWnsPdssWul++ecmfMPKZTxF0Masw2XGhj7iW9WVUQLyCH1svw8ltuzu9pwu1keDMLGEOaO1WI
NgBPD11+RtJH/YmM99UXvUsHrgJinWZRZ+Tu4d07Mz8ccNUghcdiwPWsEg5C0C1aCKfFqfiswUhX
poiTCSqQCuOCo4hDvNLYo9FGyTYKTkAq5p0Y55/MNNuzVrBGLM2dKoN7Sm/wT1/c3XLuLt35ASSf
0m88GNsfu/8ZzmR/5vvcZltP+UtfDeM2iLi2zwY4h1O4epTvzOkSuWWhy6/5VVG5fh+MVyx1MbTj
HxruvsAa3IJpXRMewsf6onMsV2xJHYRjedTdC+bt4pBLQlE5aXqdakvpJ2vCpy7tE8w19SbGmgLk
6zOZwWEOOd8IqS3t5FNyvix9bUE/pqmyUCGVnYe/pd6T8fzVOJ6nItPdRIWljvTriFkBihWjwpjF
GV4KWbGB6WKJjhAt8ExrytD4BtB6niptAkiZYZ5bhas9+jJYgzwXqzccEZLAwJ4uNbdYZfqpWIZP
co+gSJJ7fRIKeAVGf/7e2/cDFC6tYnSgclTWpfDSKksBKMhWhOyRN/6dUfH+bAEpeOvrC9R2RBTf
bB4KyvQIzBhAbQtGnQhmxzOXWvw/h3yyrTRn7/PIQbX6HFUdCf+oiYZmM6qIZtDsQTEtwzmR/Gdb
bzeEIsgwUVvTKt5Ee8R3rgvsSxPoWHuobKr3EggxRuiNJdUsaxPXZVJV5KkYRTLEq69+js8P+4i/
oclygb1r83lCWIK7L20AbNdkTgrX4bIy+ZseihXtt8bvqfBCUep9cSQQ8G9nwzZhMhM8BcUl0Tox
t1N7YcakdogAf+BTeX3OClsBSTqd/LJN+28cfVkhwKfN1NpkufxjkjdwfmektGct3+SKA0h+p4fX
fUhHG9C4zgLbIfmdHslxllUbcBXSZFjvDw4J5gVlolvHs4wQ33WYyX+gdc7J8QNk7OOx9S3XjS4M
ZdnGa/8vKK9O+yl+R25gq8Hv1eahzMj5KVcB3DY1d++bl8SJfRk3++gB88ggXEbQ7LSktOnx/8EP
mwjrV8TZlNOiHndPeBcL7Ueu5KvlJ1De7mlz0D746vyTk+2fMQYVAYRdMP4L9a082ltHSe3Zrovm
pdzI9s2hrNWTueIkw1ziclSroaY99UBr9gwayuA56elNVoERe5azyWJ6V0E5RTPoUOtdJQbnHeij
zGE+kIUAT9HOQ3phPZmzqhG4w2JqiF3nj198n/oc6ENLJZWe4WZ5JZCCLKTgfehJPfIySGKNi7TD
XOnhIdrAvSopLT0ev1ld+TWgdHCCFDd95UnSPplCiRxb9A/12NEK/Zoa53kTsVllwexixHmxY/0+
kW5M7hMldt2I/TmJK8FojccIRRvtXaSp3qwbuJYcl0HqvrIUYHPHD3NTm1DeKHWzDl/sK54InUZj
6sFBOwCIs0ZFNaQyqSU9VrSgYU/axqwmi4T+fxUQM4nu72ISAfmOZtocWVX/ypDeylQQVbq3xxEJ
HarTKRqmmRCJ5w2U6pxr3DYNm74tNIlOLc8kSfkl/hGhx0s87YrgnL61bG4QZuZFBnEJKxlolpLy
LzyLvbOL8wMelys4g98NCNQWlomp+VMG+MAUKqhj+HuQZo7wWXPutfL/n8Jj4k+r4YqFbeze+Eq+
0sTM/QUehzLMzG+jM9Gx2QRSgW+/0A3j3n1bYkMgaLkXruiox71m/TXUmQd1XW9eQIjo8xrTncjQ
f5V+RnEpwW70hTsUSfzbL0wPBhT68OJDK/YDLVkrs34t70NI35H66uYx91DtL+BfChs/hGPNIrUJ
adJPYdZrqjp6OKB6Gtx9Sv+7291aRkQFJ8aX5UIfqun14VJgQ+d1GKCFrAQa2m91J4dY9vXgSCQW
CXw9tr1t9JB2OaYlzKb3RkxztkLqWchiqH2Hy27aHFkjeb9Q9Xr5rk9Ya5LkrA2xaRfvEw9ssKIN
acyFA08gbX31DPjMGIMm2iWAFuOa9ent8vV7anOlXjx+oDAm1IOE4YWC1ZnVJWAqHXyEHzzMg4k/
4Q2wRWXxS/cIyz0yQxO8zMIJ8ThGWB4igw23XPxSNCF5kN8/hJ1Ej3CGVakTd+yr4voyOrvgzmTF
cN5iD+m55mPEDMpFhMfiVD6a/ecQTAkUzlGTQfedcgunGO60k9Tbnv5EnKYbM1EoKTul27V+qIj3
RUMYtCOJ2W6j62/tRJ1gyuhVnxqUs1aBkBpW/g9k1K4bZLnPLwyVWEs5+3v4+HbZYmE+4LAS2soE
R36sOHYoFuMLlf608hUVTyQKrt5Eh3sitQU0Kp1cpWc5oWOSBeMGdr8mxJ9CY9nL0DqSrG3yR6NL
0e616BF/DklJ5R1JAov7YbJBOz8Iv8qIl1SURanIqPNWkAzAuOFsYsHDQUqKv9bK/2NIKmsY36y3
cflFNVXzIXKenQPs/ApXDliKiWH4vxLPFhJQr1aLKxwL+/uQt3JSmxNMz3ar5rkzqyN5a7hJ//GJ
C3zspegduCoPCzEFPJL5a2idkJVM/hdPESDwkmh7IYQZp/m85HbnFvZsU3CXItg8A1lIf43rfNu4
4gPFtmy74K+NptNh1374R/0aU1aL1aw9B9zN09cDB+iv8ECI7G9UqdSZ4lFMkPFpPNxrwFVZOW8H
jQVNDp2Opjp9Gd4PZhEtw1+P47Laqmz60skkeqT2rjTZTiPiwjNrtPZbzlH0vbTQpAZZrqEKLnTg
qTFvB7vBuVFMhtnvkfv5z2CtHYoBt6ifzO5/I+a63H5PLY2cZzytPLPmHkHDp4j1yGYNEpIEPg2p
aoTFqbTP1ZYEKTK1hrT8euDJGJADTNtA3WFDa1TCcD29RPGJhGsfy609kFQtkVfNaeVFoZQkngei
OYjssPONtUhGt3E4R/ek2igfRHeDjBhC3ElruA8DfW5Ev4+ZZelv5Roz90NUtPDAe15WJ2lr0Tey
LP0ngSCHfWhlYta20Gy9udL2I6Mu4lVWSmOVhD4yHsjCGiU7WweO101DSZ3CVQ/btTi06YK25blY
ikiNg9JRwn+n6G9BZzI+gyn7J06Thv7yk1tHqJvZED/pyabdvXrjJ/RwYNjm7rSntMcWQJIPRZ+3
uaGVS33H98Kp6IQ753jGW78dbplf5/ScbBCqDurGLPyYtXYpfpoCpvyExnyeuajdf2cmRc3JZf7K
n4GcZWB+nBiVUkzNELSXkccPshnXtcMGiJdtS579VA7qPsnoSApPCSq4703B8ScxCAokEcZibqEK
BYdKcdRDZncPdtRBAT3RZZbrFaHX6VkvgFnF2ZEI9cVweqsaH6U4l4x7ghYqUYNr0qt2rj0U34f9
X/16zMGGavM8iErfQpbdhh23hXr06P81GJdSEtaVxN/Sud09jjbdRIgNUi7hbFnyakFpACaiRDvd
OLwDzu/yvm+tr63C7N9jMoKclNb4M7wYvkLtN8T3DPKR2KQojmP16xzvHIR5SzuNnkZxvMP1hQy9
BtPYRr1yi8ptFN+68i4X3XvGqbzWPp2mTmpczqUFvdmRXpIHoisGry74fS0WawLjBE2huKuP68GN
dw7LWXhNCrVxkVjo1BaH4qRbsLyve2hx2QyWLMwmJq6IrK3CxezWynNQpv9J8IdXjVpBAAeKrLoX
OuRowI0eJYLV5Kv9wSXf4S+uuub0PIS+U5lp8tLKUqFwvOho7sxVm0rC90gGiHLRsUvqIgmJHTnm
VoMmYi8+POEQ5FAb3pwqVt5A5V0U/GKgfHcxP+VbV6YInOzuKtn3KnmDxkRaTDRfr1qG0K8uws0x
NJ2tZa2zirzM2HvFUty1AmxxABWvcn/vG7H5KoeqwueIrHqlnVk/8p9PfVer6691e6e1X5ESB68S
+/ARuo1IGB+kTtlPeoqxsH0fCvA8D7aEKqGoQhWqJqA0gqy2cTJID5KOKeM9/bM7oFFaKMrn6NPk
9kwcrUm3vpl17LjgjUuHlmyDrGpuXv6nAe1+6a8NmL3I91S6noSSoh000D0LtWRGr2FEYFfXZA4s
RxIbZfAOIyktill0ONnKiqAtgqj75bt+8uZSkVxaudU7DHrZVEnzDnjbbSijUaYZMrdMFzKkwehC
fjmVmR8bYcERxi/Ke805u1W+mLDLZm7XqMn/HiVB7VzlDEZRn/lV/pn6Ec5puiG0bFSR/WQz3PyV
KxJcGlm3EyEFPLhJXqL/xWbUDLHXSgo5302oMgX6OjEpCem0xl23RxwtEaIyJrNfbnSXV2aqdx3G
BjXnbFFR9kle2wYjiPcFyBa3gVudkinWvAHuST0+BYViBL/HoGatVis7JZ4gOetVoAku8TvR9OSb
4wGPGW0hiJqC0P7J6opm4CCpvP/BjypksyCZWf/vKvQNPVnIbG7yX/u+FF0t2sftwQQ4VT9IMV7E
40c0WYH2r0u6o7may8uSx/TPHZyG1YCltsgRDKPAGJkbtE48kEb6t6LYS7WXEe3sa2JTtpYPbiE/
NswM4i9XUCb9/wGwVZo4zMl1AxWoCaHKjXr9l0MbQRTy8W89XguNAi1ZfBpSjtWG7kpkbVt7609q
q7RdA6WQFgZr8S9mVulea70hRk2KHjfNpVASbP8gNyJjJBr58OszdjU0VkWFBaNTAPGmLkWpe0Yz
A0Uk5NI5sTTbeM4Vdwbe3C53hk3bHM+iCQ4BS3J88m0MH3v7D0/SqtsHBptebIRsBrWltL7nbL9O
OfvlSQdjTg+RQh9SIUXLAvHg1jSYSMTimcwx1OVXbtLV2ljjCzVOd7js7w5DpIyIvn9EhRjBRsk0
wDOCK65ghLIMI8tMd+MAOb3PIofJ/ed3YyCKcKJY9/P+KkFgSUzLhLi6n26E/5B4hVyf9vGgzHA8
8n1/G8P7Zyd+j/lePtfqs02qaif5vv1Rgj3I6cn5/vG2iIFN4hkwf7nadeEPGBoDdV6H+rxG0tT+
CvPquqnkoFuLI0KVdD9loFe9w3cRlNiICQSRd/PoPzvWUluHVkrSjID3TDjiDtLgDjdiYXwDOYBe
CGmJAEDCcaNUAYjOFzNgzQkd0kJgcZemI8yQWbGzc6NKQZ0gixcTaJEfFeKWrFzqou7jKcbq9DwP
eSOKpv5FuDqnhelrsCFTzrSqHR94y4Z1z603XnMK57FJLJo1yed4r42vTmnDDPQQwQQZ2HB2AX5e
FaDfg/ZUEzNzGAFJNyqnQaodPgHUKtIC7G+JtlwYQXwisrIF4yn+0LyqYP/TOzV62qGqux4PFpJs
74TbR9Mw/xb+9HnOQ+p8s5Ym1yTctcXgdODSE/Bfb93n4MZqy3ZYezvRevRL2OkeCImDMoJ65Ucp
6Rbh7I+JChVf16T/QpR5B0CxtkQ+PGzvbonfJSZQ/liLKRUkFCEFKbuE1QENwB450Swk0Q0PcUIT
VDlF7py5XpY98pOka1tXYWSFhF22Tp5NplIbRddM1jGbw7g3xQwSUhvBMPZwI9qOf/Pznh6B07Qy
9+RpxZ0BvT3dNhxQlKuJLrpszRVJgsbHQX5lwaE/Rrnb5l5WFbtL4TsEa9nznjVh2f2D1kWPmDtk
vCIgTlLQgPx5IGUzFtOtod1zOzSoS86gtCJO94EyZrWRlaElsqviZcSS+dg3b4kxfNQbBcPLxbXK
Kkoh+cwNOeyJYRDiOGDvvVC88XiDbRXhApU5Fa5XJi9SsKTmCxeRLC5TmGw6H2SMh6MTC4aHnPMQ
ZQIKzEzyFxgdsEmrJhw0apRG+/uCgIBfQz3nc6eXw3jSvdn5vF/+z3lZi4kHHkn7ZOMKTAyRW/UI
jr/0/sQOh0qmcEPsSRCYNJOYI6uytNUiziS6ok7wVZLRhk6GEWJAvwEKcavQhsfAkqYDJHjTp9vL
X9SriMiHw2ZaOBBxBmTmQnhOqn6Mr8ooOEEqUjoPeCPVc5xaCFHDiy0vU5wDLxTh2JK9Fe07f0jk
FeA644L5mSyGEWarN/YNL9p7YYifSe86qzUMMKfE6r0Mugk5DWdnWLzb82yTzgngkNxlHbCMLjby
gxVmpFxHIt2uZI2eulbHEc4lhI4ZuYdTvOd4EiMlL0kjS4NHSdJpfTkaSJlEyAeLw3DqFPVHYvTQ
Dy/hxdZVAR5vOKTPwfBkDT/+AUAYtdiM1/kpM80uW/+UhPFdvLrfVw+VykH5qOIkMsp7dyYzEpGD
SvmfxZuYtuekXxB2PPARu8MUB4wfAvrhiTqaQ+HSX95FhjrKaxblbVNuiAwFrYJCgxeku3+zN2GD
YcrSGrltqlGeDVtjBaB+2Fg/sm/eiltCbXdVJ11ZXYT38NUtCRvsnarofhefzAJKm028zBdO8U7Q
oIxD1D523lgLL1iw7rD4QycCIWM6N5IWaxa6wNMFtVujdFPcJ6CoBKtEo/8Yl0BcqSmyR2Ua76uB
iVp9LbrJnvhk2qYTTNXccJ1vLvvvZS2q4JNvrbtyc5+zJrE6L6ucGYRCauz/WFZEMfVUXJnCN5uw
wjGFaisYmcufJ8KZggOqxO7M0IQvg5bXbPiRpLoHrq4LpfDnfeQWT6zpDQ0TrDB4NR3wMh34UrCJ
8eFzU8cfc9uJUaKvOxSmaCZB/T1c0nLGfi3ENJos8Jw51fcQGbmpTLovMCk8roXqf/r/KNNlFct/
zWxuTP+MnATRXtWWaNu/q6qPXAtu1JXNM8J7sim7/cO4tBtPErDxayKtqQ6CUWYHeuQEFkEftQD6
PHqTH4SXQckOmmgb2ItvPSJdpL4HNnjkD9X5zCvfvoME8GKO/swFwflcMPyaXw5aWh7W9l727dEC
zY6ipIop7qtyGBeG1bn6WLNhX/NfHiDX0FrKPAmsiTq0NIzge2d3BTW36y8onm14JBWQHGymJArU
iV0rm9CMo4YotQAEoEWJjOJOcTNyzaaOSxJckc2AbiWnUJ/oLkHDvJWKyZiy0gUpghchlnnL4BQ2
0JcbK0FGaIpaBuFiajZy5h8dwbPnuE3JrS1vSQVNtRJD06vIshk9fvYtvUgqU95VZpTO2XrpkG0N
2UzoHFZn9ydq0Qq7k46n3hU9MeJydkkl2WrwXpiM7Ib2EmfmpSVF9CaJrhkBrbppVeMNP0UQ2DiK
/IgSv+wptmvVO8mNQmRzCUogU4VBU+FI6zDPr2QexApaZbkg86SPPuZ3goag4LNnnfgaY788pJIs
WgEbLfeFmX4m4IsyqlhOh7uIbfOmRkMSB0AYksaMQUamIhT53kz5AZ31+TALZOfZKDxopY7N6yh9
/VFvTUNDcUxvk2x8zz6sRs/1eH2Pod/FBEv2i9zEc23A4aeslBKm51RbnvROtpl2CCbcmMOOTI+8
LfLPhm3aWs1Y41u6t4nJg9d5aRLa4COzW7sEka1Eded2p30E0wWEEP7GQ27rnba+1BlOF+Bg0fSk
06XqkkyvmABzRHXwXSDCOINoUQMJ5F2C1P1Gatj9CLH+KSJFo8lN/5q2d/dQ9HmkJ6ls8ZRRyalH
38gVglZRXZL8RIUn4OTHC1BEzseeDLsJ2G+e/R2349EQvdonPn/gYEvLil6WQwV4/DcvUjxEniLJ
bnnZa18hNgFq0yOYTvMFpLtfBdzCNxuOYcptHHxoLf3RJ2QHrZMqrQy0AdcYaRE6TveZwmeCTiR8
VPCYeJobMs5cD/XyBKXur4TUalioWCdVYZfhj6RxBxpKAfI5ZJh4J4ctuj1DKx1bOF/Ut9B5DSFB
wKD5V9tw+GLc0uDchdZmVtmOOtcQvYGn+7d1amVS83lq5yOqUO1bGox/RHYAN7Xo6WO6sNo4M3s6
nWXrq85AkwMf5NMrZmz06b5IBBmj8ldb0ofH93bbyuVDDEnvnPD5Izc9Xt2vAe/kCdrK8xTZS9Qt
6cktJqvYiBfzIG9XqbB4Wk2i1h7+5TJXpV078iuBSTCCtsovLoh+a2/WUCFZPCbVHIc4mULAUgBH
pZA8A6pxAxK2hNcVyrhxSU4cfJWM2DuR6R1AZ3+86s1iG8mHDVRIZXYipc75iqkaHr79V7yEDlU7
JTthFUHvSjDiIT4tJR8k7ExxMXSNaquzsSPNKjlcuT2ASIUe5ecN6KFpe7JHyITzEXFbbOIw6J5f
5WEgaHtbVvVauNF3UUy3VAIso60wI7TWTXSb1URsPLrBiPymqmLyiCh0yzoRNST7LgDdPOwfYgZo
RYb9n4sEzE44JwetkdOyzOpr/mjVP4anCuhLoCSezU8Ex92ToqkIoFqqH/G1usIFgjEvrc5zK2Hz
wucoVg8v+AX3dwqvMz9f9uIMlJl2RibWWi36ZTn2CUECYCgoQNZCG6mvxn/P/9YcYoit0R9yc7rz
/kGsUgLxg2yGORckltW4BY82PG5r8+bhrXkGLNHHHspKCSWJLyUGVxRbWPfFADqr20VPjmTUDDFH
xrsIFynp4ECuZpQskeRh2P47HhCzaAf73snev2KKbySyfd3SE4c2vk+/txKKlzYuhTytz5ksoZ29
5WXcwmqueHMwE28Z/xQPUFin6Y0uJLvdmXCupnGnCaDq0trrl37Zl2lX3yty+72XPyQ5D7lrx7LT
jxXw1SSrEAcR3yuonOmatpdUD8fkdQSFU0PWXjr9vd55X+vZmWlzNAjFIKo1nr0bw9U/ChMsWiJy
UoR4hUMp6bbgPth56gfPiAqQY4/Nn52woTGbCwcydSHVDXnOQuUaq7tADQorTcOC1PLM3vBKiip+
9lsAaze3th9/wHeSOOKQoKZuvngHAt5uJvrwxMbESX9lT1eQPAoKE6tB6CTmm0dFDwC3VDEeQsqR
9RRh2np91j2VgzNuypa+rP60mrdPDWEllrrkjl4KgCswtEGIKMJcrkxPIcjz/WKuIBFjQFXabpnW
RYb6wxbJaxj3Dj0M9SaRghAPLlWrRRFsE7Z86FaN/Fzpzv3wzR5/6gdOXzm/TyYrStO7LK7XlytP
i1BCMh5CFZJT2zbyJOPnEklBf8BihL0CSH6xkPl+6B3iFUPtnYbWQ813PMhnCxnuq8RaH4HN2hlR
DITjCqiZfGQYmW0xuzCmqXsK28S3J1KMF3J6A+zL6lRrpLhg5EDEg39Q0V1ksLV+8vSAufxW0hNT
PerHhBhX2BDJPQOwLjoZYMnTw4gzk4+yhe8iIF5Ea9qS+Avk9k+BWIIfub/NiOFCEGfpe/uip/Ia
/b8ZPZfdVBB6nTfdYpmTrMSkT6J1YvTt3SjdfOvbPA150gVwdV8Gh0f2c4ZY5YoghHeDs+ocdzc0
RwP0/5InWlkv+M7CTEpRZrGNXk46ojZRhuWea9mexjpQ1d8h3PEf1Sw3qXO5WthN2CeBbdfAnayy
FgAZ+VfEP8aYaWq7xUj8O1ewqig2XRk1+aKbcCql5MG8DBa0u3ORgko6TwtJviE5I1DdKEBd+2vb
mJe9x95hwSS6zj737NxQ1SkaESdAgDGwlPWKq84w+RzKh9u1eVbTehFitqZsxIwpZAATGs78mdqk
cD7BgU3OSgRUNPskoFCn+8W/uZ/Mq+sLpJ6/unG84C45rKEXgfQSAU8E8+rREEHSH6cPozUPHN7P
5HUJ8Sz4lNUmKNKYEQAo2AJ+Mf735FteaA4KjvY4yoAT8bXAoa0QobcFQaIB5o/vD7ejqgzRfxcL
hkCa6H6p+GCL+JkXwEoXs0AnrLih1phE9dkoH9r9Mwx1MtyIW9DT+uZ/6M6ITLUQX/6+9CxtPakH
X9zjTwA/+awuZrVM3r7WfeAqa7a5QZvGEFXQ7HIcXiCN5yhnZsiblXZhKrZLOSbm5Sd5oawPzit5
t1XL8+8sjaSxCFT5DDE+oCZtI5pX++ihMwclP0RVs0mavS4glcGSIpsjIffuEZ2AbSY3VzU65wMb
BWh9UWC6pkmk9xsGtaVD9YRHZ1ctWO5X6FLEOJ575YU4p/NsWzKyz9P9KJbOPj6CF15KVIGiPUoz
EWAwI9dM7tSbBDGRsOyNFBuC3nb7oPTb3gxA1BUIEoJkQNGOGtKdc66ZnAvUnecUZmED3GsTd0wR
s5N+nwutERjz9CkA25OKSlTy4rav8PhVuM2nZ7bb2DKW4agBjaHTdeUJLc2wEyMS4DnyuN2J+vHI
/62O/QEKHVcKFnJf6N3ACbWgFhO8jdm5MeMAny5yxyUpZCLXCBPNEVyzUyR+dQA4fOKX4Sz90O+X
fb3rDcP/vADC/AEg3Oo0Vlp3V5s7ABFiKLF2nieAuGNWZP0pxYvSDdHvob782ZBV8n4IMVxw9qJW
vaQGDlvtBPMkfs+pmHageOJQnEsFTSWWXgvb1lrJMBXxnrSA2xJir9A5TE7LLa5kZ+fKNFPooHSC
bJtczNdD/gx2CFNlqR1tSMG6WbTogJKGkgiMIn/6cwBkik6wfiHtE7NYOdW4vvFle/QMrl0N2363
8/GGqcuOlVBZyeKYPB5+8H4lumm1E4tAaNG2towWzvMxv8OapLw+Z89F/88qkR9G0mNld4FaBhrH
vXPOqhNHNCgBRGxGbjbjIUm6z7wE7un70d8oP+IqnK17evPXOLqVE9fISI60mLny5qI/D5NF/ETB
foNYvKhK5Sg4xEZhkeOyVXW3F7rjQwjPps/b96MuRidpEVY0o/Ajwbcw/n+k0twAFveVbCCw7aKY
LcVazH+t5gkuKRPyInE6qg/+Es8VlO0j19fpMmcO/qIy5Q3BzkbheFYjy8H4rOB+dr2AgfXu6XYd
nadsF2RfwdAPYAbsqXr0mOdqnIxh3Ga8C68e+zdh50+mrPVSG+qvb7Cn8MftPI0R9hmM5WpV7VGO
CoT0v/P2xw1TVCMJvD3V9hSLXyG1whZOTT8heyZg17sqg/ia6/N4zr4ywXXtLt+zq0aailRchD5i
WwoPLnQ67D/qSzuLqxClyMfcIzqcAzI0RNpw0IIV8XGfO2r9+Pp7RDPWrtGHjQisV7o3wp5rKm3u
jDNZEnehzOTGWygiS5Xed1Oa4okizoopuFwH1y7zziSMyCaNXgd5Ud/uBDSYe138WYTq8vZfjDxH
oAytGPsQJJsPJ9sBa2FIb6O7zil4C35yD8kKVvv86IoEgcdzYknrbW82CWFtZXvZXa8oLrYLDbr8
ms2xwPgAoAHzHCPHCLXZvr9Axmw9Ua5NJRhZ4xkfojmo9rhEiz4GXcvJtkRH6a1AcM05kBuYXaHm
Flerm3N2xdG1+ChW6CBYByFDXb090fGLwJgAztghGlpVrG5yLhjgFrtcAe8aAJZ3xEdxlqwZJnkE
nqSc2kYzK2zzFtZmLSf2GlMmjezJfdwjMyNaT21CqmnngrIDRRFlyXSUG5Po37sCWO5jwOqZAMCZ
ZLP1RWz4dwSQtEvznkzqIuOt6rsalqJiO/gEUohNjeUuLPLJrEyOjJ5bDGo3re8LbMl8gpgcsXx9
p7U8bIGspEOss5gtdW206XBR+QvhotOVVsqyjQnvlIc9Ehn2YQIvw+mJgP4BWpbXnqtU8UW6DFxO
PPFgpdsMyCZjIDtzVOwxxY5VWER3BHMsyzMeEX/AuQtBOtj9D/vyGsRYj9eKiCi12PIaPUTjGgNp
Zf9pWFRWqUGncFFGCdMqCWTVq7h0O8MV4E3wkOkNoYBgvHKn14KSh5p6+YBj7X7fqHsEO0leRTIX
COvTeGqUQkoZNSx1HDW7TPJ9PtKLCdqXewoAZPo2PvHnlkGgbVyVxb/TKrkL7rLmy2azGFo5eDEQ
PAbBDdwZOFdOF7S3w1+JOm+dvzYw27R9pfxCoRkZND+UWc/YPi9pbYUwY509k2nQUXzJ5zWccgTj
N9VohJY/iNtQSYweOs6RCRdJFbD7kE/ticKTfgkr5rtIiDxvYrUKx/06AURfA7ExKE3We+L0rQmF
Q/fECMamV6JMKq9QuAVzGWueftt7NuVwMzD8cv/0GrvMRN0h18lNNHTvLutyN+IfHYQpcPG+PNiG
kyxlHKYxHeeOBGRalwpKuOTQ1Dpktxw17jWV4Grx4ehbX935/ykAXMPafZoXkgwQNcg3gygPn4y2
kfUbTCj47Fvc4XfJvvPjB8UF0DwZIb8QygbXaPPF0Z6a6BTNXLfjrfrYA1eTTbviIvwze2zDIBRz
laRJeItByBoeKNi52ebnS9A5e4+U+D82WTbBkbFSvmdM5BKYbU7I+Df6pCmOMWjm/zB4dpjhEkQd
PKnrwBcYi/NdinlXc1Q72CJ7J5ZOIWSCym6nuprwYm3XIJEcRbhhuH3xbNLT8pjTOHRR51dlzg4P
//XbpRxSv3zQqSzrB/qKRjzQ+x4xgFYHGnxbjMPZ0hdVsRJVuDeDwL9O7ZQyyZrKp2ta0bxUosWE
43FS7uQno33VoJNuN30SBr1hIDZkRsVMoA9R2Kwj7oUGyAdt/Lt0e+KAghHH0T09SUC0MHYu9vko
JUUBLOEl8QsQ8IY6fhqMFMNakY3k4lGfhe3jZu4I/U0Pa1IvqEhb8Wcn2sezI6/NeZSJWUKgXNN3
zjMBdNEjUHY7gbFoeX/A5OlVYqSFqRAcMycyaG3lHNRnnjlNAGnBlyRU9Mt/HJh2vf+v2IWs/DHH
u+3pRV1820GyG9bzDiPGdNcEcHb0/OTAAHrDyk/uG5k2v5qgfj36SkZ+8B3brGx6jVbCoGR/ntCm
d6IwnlP3xNYrdy2nSwCxHV7Ur1RslNnavbw4a17rAsd8ibC2d94ZfPNbdYKvAKA/rpH7wqQYPYk1
mf8HP1ficBtV7gS7M3wq8abQNSAg5GfR4CR75bR/j1wyedwvmJKfz0gIaR+/k1YyoUjtt0uyYOxS
1erjP4H3cxOgwvdfVJuF4rmnFPJwXSQdU105I/5whtVw1fqpgFfRA/s+JGkEo0LthFjOITcGVks8
fdlgx28juV1A1fRAY4kGHB0uXkHLxPz+h/68PW4sZId15LKpn0P6/FSVZADn3vi8XW6xTqAMC16l
ouYQ3iPXGx+MseLFDr6/mhqbY0YclV+U2VB60Z3TxiPhgiCtyfOKerqD2+dAjIAGbalUxFLa7u4I
q16mGVScZWCWLztYtKtQBBW7tOzqez9m1cwbwU3AiTCq7USRoknVZ5hARvcd3hWMj+JJ6mVKWa7t
m8ey97N4Puw8HmTHeZq/Z9vw+mQIAL9N5hvk47ItraV21V7JhPIk1RUXkFJJVPFN5BmNR35VJGNT
3UmakJ0QfXvMd7IKH1ux7v2ClTYHVb+5pNjcqwqsuktw78/ifGro9DRjg77Y3HQwROf2YAunEnkW
nArghTd+YgR6LiAMDJN5Fqajw+EvJzu0uahfpBeD+m8dnWzX92AkHBvcCgtLSlkEZ0b22ML9tTHh
asWpuoHqh+b0/0tF9zSgTl+xxS/uIG9mN6ZtI5j8U2ICy/++GBAo0GGXFF55Rd9q+jVS/S7yBtg9
QVYZkg+Zrs4LrPqF7NETU9YDILi9zN34VtwiXC5tT/JlhmBph5fz2XoudC6N2ow+U9a9b7pRtOAh
NKFbTKp9poBGUASp6n5Q65NzQlLbQMSTDEK15Cwhz5JbNQtPpXwZuKBf1QMo5T8Zzib8XWMNyxoe
7V5f4B07uP/p7a/3UbKnWk/0TmkhgsQV/zmY/cxBNxpgiVGvWPpQcZWH1GRyRZgat8hIuI01VxBy
KNwB1tY4Ru931c6wpq66Y6jwjezoVXZIlIaB6xIBdhJXZiXd3UYcUdstWblunqHY1qLgpnEcLeVx
3tj312PYeVy0QPjknClqZQyyHf6quPFqal/diuq61PC1XxCOggZzMFrSW4awiQppPsb6tQvUS+hE
LWeZgGudih/U/TtEjhod/nAPU7Px+dRAXweqrddF6BfLsCjHvUIW5TZGmSLLLi92BouJOJbW7uc3
pu/HqyU+mnPwWx+bhQdCuE0WK/nBLl+vrAEsq6y5OGdcc1vYIeThkT8chjOWEoAX1i/mL3ut44ds
ZB1w51MwtwRhLSb+Zmb0MorZTK4eTxraWvricSAMqM4H5KFPgOvVRuJHbrRb9xmtdlBmo/CtiE+c
o6Qx5zsqSG8bTK1kF5LqaRkAmeVXPlvCKZOQSt6DVYN2KcstHhJbOkl368A7X1+M2dUXtTTrT5LF
Em5e8gAkZ5Q1aKvbl/qJynKKhJ26iPbNUvix3K9gOburfPJ09FU8nFNZMCj1opN1b1TOypvEg5cm
oif7spipBcN+9TDgbyEr2BKj67sosoD3Cp4W9JugAbOCVs9Me2F3F9EJsRljiz3EdCTZSDiXoOBa
X7agdXUWqOlMCuwf+ZsVdwzHgwSUfrGF8l8Z5TjeIUXF/M0TPyfsL7WD4VSH4E/fQqixNEONSifF
D1XujDHJKhzVAvUCGlb2nr7yk/ghnW3G2s0/+TkOlJRr6xXJ90uCLylH3j2hH84WSsUEB76V9cXJ
Wv1Y+176AIFkHjATYlrjzRbGAFZ6VdN04qHI3NXHP0uoNVNcq1Gkm3Gw3J2UNP06HFeWUg9+df8Q
fDeGTSLB20eYztdIxw8PgnXaBGmjbjMqf/2ej5OK/PKemLDdRRi9k099cy194fKlzko5+zBTIgoj
ZIv8mxXdtfv5cGeq5hJTeaEoYD0u0yfpvXAa1nCFpUuNoJiDHSMEc+i60OK8K/P/1Tj1nw5onkgv
kUzSmxHo43iKhOMr89XkxhjmnfqjEVxF2uPslIxosSC5+WFmQrynzCgVx+eSB1wcabYuR4+Jhp6S
LW5Lw3ZXdbl+OitwSu9pCjaBMIMB/rzarcj28Wj4wuS2cfHgeIUkzivEpOzZCHdIfaDl8JqIYY4q
+UG1qhk4dXRguTpgUKH1b+iOUGQEZ3uv6AUO1D+4aS7GxWLF/xS9C6Cw9YrqldIYyNBNywcv1isR
aezCNqvmKrYyfPgR2wTVhj5Ff9mukX0wQY/yBuhaKMMaGvZiF+d/ceDzd1X0vlHv0qWXhQzsH+cg
2sxgLj35FO/Ko+J75Smjt44VWbi8UCQHLYz72rkO5dMN1sMgVqoQ96FVs72XT4z6K6GVVWaSIKTF
TYPAHvSW0zbwSJdsllmkdXd+Wq5hNHWgfckGEf5caNORAB6WKGGSrkBgDi0UI049SzTHzoniEWSs
gtKOJtPrUREUorow3bfdvXM5B7xauNqsdH0CcF5NKevva7AUoxOyRtpHWYz4kRTzFTbddVNLWMmn
UEbz9hFEoAD/pwu7Ludlh4AfN+AQYDwDKSDwZrqAYsP2vI/1LOvkoCP2bE2McJlxPhbVPt4jxshM
gatBUJRTq95fOztZFqEO6+r2vD1RM9OAyqE/S3UnETmIXo/j7W95uIxgn9ZZwlkSFN/rILGs5AQN
AfzOwWSlmTk30ODdaF69GWQk7jxrjTdYl+JhZKbmV2W4qzk0QxjXX7C90HrCN8/70yEp1JVKCZwj
7o3B92g+M6XclZEymzUz3m+sQ5GXm2s74MwkE3MbiDcRFOynq6l7f5Q05aEtbZ2dnE7WJSLgn4Z7
8tGvlL/HJsf/9DTnBc8j2JDv6v+CynfKdejU3IE7+QXtFX5bTUqx4WhBJ7xEnNi3EVI3YPqcDsbY
4Yb8/CbLnJi0d+nKo5eEfVhnkDZUP2jJdaQ9KQoCznW6XqdKVFDRYGVrQXH3Eu2vibHieSMDzZRI
YmVc5orW2PmSKuuTfqKDXAS9MOZpi6UNzNN5ZmZkrjOQP6m6ItpTv2fdWcTGSAKNy37sTJoOXiu+
W1UAHbFuGfjXtbU4G7uQs+175A9K410stGlrysmA3hylOvrsgk+oOseJep1c7/VuyLCtwXs2gM+z
byE7SUJqWyHXsoSoqgYt64kJ88OBF+8oI3bqmUsrKRh4WKixxxAWS/r1KjTFQTu/jFpV3cOPLFOF
SVka7d+yFIONweDV9TU4GBmPAHX2Sfkpf4I//RfKsuu+nJjBp+62AChaPp8K7FGiizoO3y9EVvjn
f5/wfZG5Qa//Ip1cyNmOd/v0nRmaIfb0GQ+pQ24Gx+LbDGEFKrU3rJl2ip/TKVOqmP/jxV73xGXX
/yjZ3PUfuCpqYsR7UHqNTKH5Y396BRxkcyAI6UF4423TT+g2t4eoTiyBKPk04R+2Ul5b0WFVs1xS
Ra5DjIbmARuRRYWKrFFrZ5eHXpN+K2s66+2DXI9fUXIbC9HzmuUa6FK0827pbVKU0kBg64kJT9WM
XlIBOI4S/kDzTrXRwTYSeISLQS618HPpm1Kb1c0V1FnHwwRmREv+qIWcohTt9hIkFxNH+Mw2X816
VMQjMdT5i2ZW4hn+09tBvC8wsp8lIZescWgTspYM0IyElLCqdit0sQtxB7wGn/0liGc/xjwoNnA0
yCEEbeOjbqLd8s7p+JFy5xjE80Q1v2Buhg4biFnRDxxlgA620Va/j/YdiZTmCyi2BI8mv/VdXnPh
hxlceVuLLYHxY+YiMNIg6OPbvg12DYa89xtx1Q36NGVzl0mHwNkSL5+PEEV8k6Qglql1iEJfrcqu
d4l2N/MpqjpiPZxn0JIwFN5MfDJjdMA9nmqVhG+YjxCCx0XWVF4aQUv4GmEzjRV9XGTcLVo0+kao
34R9MQDn8in9zPK7KuyqQKuc4lfN20ZMY0EG/1dMIBYN9PhJaucnLW1vt9upEHT++4MhUG3C0ah5
2mxzOJt0968yq50W+ABKE9VOKoF2C0bWtRClhdAGMctMtkqBkSc4XMEu+CzkAJCv/3G5p4L3IVtk
7G3U31B6RgtO2AVxAf88T6piFohYeDeRmQV7JEIlg3r2ShcDDD/R4dc7dn2eU9wsGt4ppSzefwkS
ukmnyWklecZxc/gRA+6pcKat+no07PwrD7eGuK94FdwEj5rDC4inN0BzhxNzmvLot8N98A1ZutqD
jK99WnRC/4rI+YwD9efGQVLxv9kaAzmF8Q7Hc5oGFJPe3LVoY4HLRtrRzv0ppbZbK+48VCvLEaAR
84n16xeSShLAdLzIL4MeLLeoHyLKECbYymvKMdL6Rl9y5aqU4vRp85U5LyGejDgfWIqbbuOtrlW2
FKhuCYEBV3YEtVPIExA0BvwdtjaiY1wsC8T3bUDLSZrYNt7ufurRlLJdXtgxbM02izwWTcdiztFO
eAeYoQPwc1NRhEoAFhF8KypluE1NOVpvwcANB4YbIWDle0qnGvq2iifZQfAS2l/86TVjTYfKmLL+
Pql9QvFmweCJID+piuvmU6b0Wr1VZAGdJ1EpTW+ZBy0+ai6rntBLyWjr2gb8gpnaLmf5pCEpYmcW
SAh6ScsZL1P3vGxvdCx+ilJyDSGE6LbG3JCVsYOCtrIfZJ8Mb0fu0ZbcrdRsjb0QIsSV4oqwRs7K
QcHqi0mezS7S7p4uhYgHaL3Y6k2Q/YgtbhnYPcQtiYf/5kh3A72IqerIGL2bfu20dYVHkBJ4I8Xs
YvdCeHtdCBQZ/EP1ADvYiCTdpNLDFHxCcnvwadMLdkuCJ2MRbhwheOJURi+IE4lGMj7ocITtT5P1
Y9KT1rf8PfF7c3XMkdHqUhrS9FqgY75/D1ojqZM1WDdxwvj3SJewQA9yuv1aNDFJ+wgLmIrJjFkA
4bKmMefCrKek59E2thHzAFQ9GIU1XRqzVedCkiwJnnOlptKQ5eRpe/8GO3D3YxAAj0WKkg0bnGzj
xT2oBsKwqcd+vw9piUT5PaRN4wsL33+fN2MtSzFRuQ1sF+uU+gXmzt+Jg5pfcydmkr8ZoTeEsw3N
oqFDosbXkpf9XYxXrE1zlR1fFEeGXGzS+t19ugK4+I/d22qsYoanZS4YPNBW7lu5eJeV/9jKkpmA
GLD2DvN0nXRTbQwW3aS/ikgfeT+1e0/Yjb6I7eLn+DKLI4AU8RCMZ2SkoETgHWD+a8UDWtZPBVxi
EllG3EpomnHHvplO/bhCsh9+IxJd5Vop12g5YSLTmEuD/X3+FJr1gbE2Kk0l1caPH+zZxWOywQNh
Ldv/SxpsOeTqZkW6FhchuJWNCgPT4Vx/R/vqKKBGgwyUiQx6f225ODTwndGBvJJObdLcDVnEDCPQ
Nl91lViQRaFm/DxpxyiePHc2yijphsJFNfTLXDbGC32q12cogYV1K9Rna34lDtxRPOJRGw+/+VCV
x8xQ81Rvg0DRSzboF01BQykp3aqNKox0iFI2UlU42EbY6lUDALal7AftSpiaBBPx3316XrWSlZW6
oVCpeTpl2rxQ+tq/Rd+kzwIML7A7O/gp+8OZ/kJmo8whIAIpC2zGhf9O38EJOjGz0BBJOMVv+SLs
NYr6IbbttJhNPzCw93immCxoXwzMBeLslnsInyMUFt+NMx1CPvqXbfJM1vjCJZ/KtPtn7SXU9Amp
nHSaLvdt501NpM9UHAOp1NQKB3ayYfz5x+tGNqZfvKBnFwjBoNjMpo/c0HIqDItoBZGo37gC7nbY
qgZaDt5eO2FM0SyfGaBnrYsvwi3+3B5D6umw+jRbCNpEycxoF3zBWxfSMeFzK49JNn0HkKuoPgOt
3qSG9WOXYugNgnisDtv+kOuv9W98wtcr+QUADZL/skcHUG3tZ7s7rEMX5Z5KzUfu508ursqM4XPU
oRyGCIpc8Zh2PN6MRgTrHnhMdHOK1larTSwDEl37XdnqgMxxYRiyoP+HJkQ3tWMd8UPmiqPn+LZR
Z3ez2pm0HC5K3cFUXNtMGf4N6lAehQkSFigYYG3e+AstJcmd0Harf0LKk+zXL920R9hwz3BwWlOq
HetY8utor/P2/oMwpB4q84vw005R40ce9sQ2vaAJaV14TrFSB9zrv/CaZB61xdbR1xr6ROKQN1Ul
SR/MtrwZDUo58nWxzMiP/E90OiIt34RdULuRSVis7hKO00cn9dm7eVqEu2zwpJCuCwuNza/tTkVh
iox3zhpB2b8/xsLlxZVbIlq3DiTShM/N4SwqLpO8QTAsA6OvqXeP5hhV/N3N7P4Afvq8GAtVW2CI
1VY+kI1NHfkoMtDZHDv/sD4dGBxFoJjmj+Mv1bQzH/K761UMStRax4RXcfX2CXPpF2Z9TmqQAISl
ywArScWAu2mUqDD7htftNZBR0Nw/rJK1kS6Cv+HGc1kTkWkGjb/nenurz1Ha5D/DFWCoJr2LEUrV
fTLpOooSfQ86mBYj9P2KywKFhn93p+4vaAa7bJtJ+HuXJQFwgEYZ1pyUWL2AtmQDfcgNj9xg6uYZ
AQ1BcTPNKMRQ1n3MZZu7cDXACLoBhAaMJPNPYvquKHUJ9l7ixajJ6tX/L2XmNV5gexklPipjzVQF
XfL78Tx0zJr8Q8kx+d998BjWvDfh6Xjfn2XDDa08NmTvATBT1iln2TWOb+Zoawvdw1+pHcwEtaRc
svMmzl9sb0Ql18KgJa73nv0l7A5yOh04+8XcaB42xh5MuX//pmpmhIsIop87a7rZTlU+mQYC405R
cEfF4Q9MsJERYLZzyMqkhYew0pT74mqr+K4aNx8WbFbOco/MNFwa6rTJDf6xU58F9/y3MV0WTJxE
NrhfZ6qlnW1TLFyCfC0Jgo7NfUt3UxYCY1rmO72kFnwJQtSEFoO0vczqi/JEp7XOOHK63TJ4siBp
sJl+nCPeqDrUW+6TRehmZ/cwRVxmxOb9drd62wGGilFaQySwtL4vHt0s1F0R4FycIOw/RDQejqIs
zf7BjkqtVF2Qv1gq9ibNJjvH6RPyiWzHBzUq7c66Rqhg0zmSZcZ6UQ/BlZv+orErYKceXaVu+TgU
E9j7dYr9Yiax7nppT+bAD9wVSsHwgX0U//WKdv5ijFYjkE2S1FiHa+KDVS1MI/SiuAv9dih/s6o/
fH6ouPXfOax+Cdrt8tzRjKXd6w8sR7KZnvnTQ8/8m5cWM+4ul3bhwdt+1yGhW5jdhDR4s7pLDIPR
0sqKy6mYwv8kYxtXFSQQCkyQcEBSSxjAl41QgU0ADCexRLvyEAMGxxnUBBs+bPUdxnL5p8JVMCFe
+qlr8HeGQS0q4DFXUYpGdN0R4Pl7agpQiGeYUx9h+L6DikpaUtDOd91V6IPFvSQWma7oUjwOdRL9
/R3+TE6biLtDpv+xs2jL5hMm58OPd4h9gSK6xkSwkQOhiihKY75n2zfy+LCOkVEjhQ3DQ42baW3Q
YT3gwvvslCqNfRlrrQXqbKBo38KRnf1SqHvfuAem838G+PdsHsITZGfGIKoqqRgqp6FKKjerLr8E
28ta1FxPzLvkvRUAFQ3zZy87zXa76azT5OokczgcH5/XpE+YSFzBaTV0oPluUSpsvJpgBxYRKV+b
YMKqmKWELE+fIEpOI5uh1o14L1GF+F04dxo0+rAdEnOgf4ZDVwP8Rfl4CPpIWEUJGB9hTTi+r/xS
9M6BMS8V1WiTvPYEK1PmYUMyQqHlTcHiONy4No7IHisfR/RwnaHs+E70Gaxh2HLgw6H5IvOrFwdv
df4hHs0D7WB8WoTCcbULQCJhQX13jNZSA8bdJihjPrla/0bCxKzBRyrLweh4aRKRqu+EHtRcN2A1
YE4fZ+/23BGZPJU80SYoinISiWx7PPDbNXzHQB8RYKRUshvQMi3hxbDeAPMmKH0UPEijDm4oS4W+
LQGdh8dpB7KMusY0GF41R3V1VoFUuPZIdsdCmrihnQdxLioahC2HWgRfoqRH2TS6FtHprgo0m/i9
Logpeq/LZhSe5iKbDiFsc3LxtttwoIhClNkcXMT8ZyRFUCnR28Vvb1/uXX5aMGN5cfwwf7ruS+hh
6QKltnfWFxb6Ozwmdsncb7JHcO10lNimtpOlK83ZGpLwZbYrWHH1Hf+7cRpzFnCulM+horLPg7yI
1ZbwanUX6cUvrRpYZ/kXKD0PLl5naj3Piq1/P7aD3bl9rszX2aJ0EcdQ+w+oqrr6D3hb1ATZByta
tilUkEBj/O8MmpKjhFg2goitvFjPhQ2jFvzxshV+sHFOhdavQe+dVxCcBL5w+MvZJkDr2f+nxvO8
hxcT7PvHgvYKhpqQA0wTv09+jGQ/eUxOvq/d1bjfpJhn2/cs8AFRDN2j11voA2JyVVh9Iu0Nv0a1
XXFzIKsZaZCUKe9vr3awdrleKeMEbIWaxzjSeK2cgSr+SoI/FkohfDIQkU1JPAc8WI4ASY/hrzkF
hpSkru4ZX7UzEgfLAenbKQ4cDNZAYv0LN3OPlUW13OsizB6qhv7HUA0wmm2DvEPaGWwKFKmY7RyX
uh9qu7LY5LGSGTrkwX6U55TDH7jv9vOJyKeYMIHQt2hJjIYu3cOBSPgq5a/EAcRLsDxuiZfeaNgG
04A9y4EUusnzSi6QXvvd4gMOONmQ99U+SzRpwZH4msctdR0ZG62Zb+cgCd/OIIpOBnPJgUk3kcBk
O+sP+mLPWsCGkWr4hEhLHuuiURVm7lmpnY/FjFizSOmAjzdrdGZhxy3TCDN92s0OOHkdP6YokKZt
EITLdfLQVLaBxBF2RP7MkY04L7PymSgQHaWRQES4BHE1RGL+FxH+TMQVXCztd9ApWT1TKcKBrZv0
tCkgG1uL294R5C77TF9cKLNDBRxW6ih0+ejMwcaSgce4ICjYJp2U2LHzx8nhIOthF8keMGl3OH4U
K/yzDnTgSKNjMwsZefddZGVEqa5JCgpd459x+er+cWAo7h1CsrLPDb+dko8dz7STCUyIDmisM8On
yWyajNICvhsIcQ9MdEpdHfrEWhTmWRCELkO3nIyXygS+VpccgGWQeUxrjjHLviz6TW7Hn0FK/tOb
3kiAgxkYXBWTUXhiYWV4/mNdKxajXopynGmJTiZcAwIy5VZoH9bPCWquWEJEW2YNkwtvOdX4y/Ew
vQx/vbGZixu109qYwgNpvwjE+jKm7LLcu/xpH1piS21gIl/UNqeJq18O0IFcmOLXJo7irK8GYal/
Naq4EWsg7iQOH0ePo90V1nx3mHRhHC3FfzuDgJuGuS67t54Ka9pSVsFO3MMMtsXMebbZhBNubdJo
50iY6tvv0bwpf6fqNxhgFfKgMGrB9auhi5b+3FVdSGeilVY8QJj+aq1atNRP4jo71WqGpFgcGjRe
MJkc8473piZPA/E8NaI12Pgic+Nvqu7FUgoa3uEWY9OPxDsEH/dchzVi8+XRCjwNl22cNsvJd0pF
FtySL1L3ifFRNZsbP9o3IkW+NZkx4ZLbxMCAQkqXI1RdC5pc0xEjhceo/cwluueppjo85kizZjQi
c60h6dxg+btZYqMrRMAZhzi5/UBt8gAQ/dvhuPaES1v4k6d9FDrxoi95EpElJJHUjaikq9oMtohE
Y0s1qwZzAfgW+o3uCbK6B/mgHAEWpfoMFQzRYGsJ50L0260mRtAtdPQO5IBL8A+vXTrHA3foE+++
FykY96L2vx/gBseiehCwVexVYTefnIdS2AvOI8XXH0f1cra0XrSvrczJJptw4X4mWxkAq2oacwYN
QYpBUzKtLiflKaC4sRbkZ2D1sNIpO3yFXX2msBTUiDKJn5r5zxwv+zM0uc/ioJI60s7PGDeLQxMo
8S9O8JI21smkMCXvysDvrhP5Cu94Kx8YVNyouN8Y1YTVKN3wpjEldxH/8qkaGkhzgD70Hf8Wkstl
5+SsFCw6/Xgy9VgOs3DQNj0RVLY5N8Izr9lRe7LdrIZ/nTMjtkP6sE4E9t/PjHr87TShBSAWxHAl
8y7oHW6HVlB4Old11CpjXmYGpMIS5vpbVdx9svhYclTuWLibkhRhfdGW/lb7SGdxRs2GEWNkGtiw
TKvcKms0jqBzBHqGoE73tIEZ7NV9KrmeBwgtWsKjRITErPPGbULD43vJPurHlW3vqexNcFzWvlQM
hkgSurL47gOlT5/gCoQg7vqunrxKAmOd4Pxl9Ih8ouhKo3qFhFecYRPpiyw/a3qLi1ldeP+L3VIV
VQUPlCAot0kq1sFbi0eZZOg8xvPfU2pwWhuvQxbXv/SNNdOuOWRHzfoP0fw++/p/yAmorh7XOCTG
soPbQJceEbS36ZyRO1yVEkDEPGryfh+dxtD1eBpqz6QGIXxM7A6o6WeNBBbo3qdv+oLDC3lqy8sX
o2y7yihKEnENcuMtXqZs3YE7eRfqYzOOo6K74RF5VTt1/U0/Q/jC4dkVqcHpCCmnA2KovRZj4YkV
6Bm5Rgce1yIinCiOPWpKW1D7e4NUNmZjDtuYyOqpncuaE37/F7JNtvOUXmK13gfptsB612HFWXlC
a2EfErQ5QyWP8DKpW3JTpsV0EZAAuE7cO0lRowIjjp4vXeB40ZjSO9jdZ2/iaSqLDTAM800uLdQP
ugTky5hltH6yfee0LIvwE8EToli1dg4aNQ+XmCE/hQuobkfTZJgmhr9jFWzfMODV3O+4bImSeVhl
6mmEf5BpbdcX39mR1pvdfjO6arn5hL4c9L8WseLGGIme/sHdUhmfD7BD63yqoGSsI3NiCIAepUak
nbys6v1U4hOgP4RhxAKvFGy1oXL7VP+NBgqLfz5u5/5UqBFfGnmiZFx+Wz1rre/t/4lPww8jqu7/
RbqVDpyY87wymkgKOMn2zC31qO+KLYjnb1186z+h8cOjD9YN0xGNl8sfq4W9xi6Yeg0qLNLnPHMB
Dx10AP0aDjlOHglFEOYwn/xoLFbEAmBylV9TSOU9rwZXe8nmVRxAh/GwWbWkwph4aUvNmRiI/joz
OSUD7yvGDSdM9XVeNukS8SRBDEE+WRvoS0jR6pXMokOqZCmqkKD3vwPvwFXGkHHaGB5OV2Zo18zM
bd+pLl9V21A6zVI0AWilUwMynNTklhcE7w0hZpTBEpnplnl8J+FGIq2b79qb6bqJLxJzmq97itjp
+LbdHkZ/4ksB8PNi6IW8tXkJE1/E8fsowu7ui0rGmyC87jzzePNjarSgLCJYmiSkw3C6By63vQua
j8dBxbGNW+oE9Vshkw7oJ0NDpAXt/28XM5phDk6Y+QMCj7kriIV68AtE870Mg+0ms898XfIm5OAm
0df5iD/8LxJf5VLCKskGFthYXOgz/uGAL6aiWyQSDbrmMKHldRfGMRuklvwQ/3G+bYVTpWFvebjh
Awj7+txJtQUFInfiTMQjSztSzfFjM399pcPl9QBKnDmW++BC5In0p12gze6X6gmh4LHuZSqbLkDL
5bCGvgJiosOWU/FOxblzT15sEo1ABF81cbuhfIXlT5umI69m5fPuNDX9tlyPf+77S+sJfBFVocgn
ACA53AZcMaYbyHeRs/fOlMS6FY5JDQDHopNaG7iCe3nOa1zzntsb3o3Wq/ad8UOVGjpwaLLainOe
Yox8L+6gUxxmGkJm0gff8G8HH96XusFkDWuCmePYUQbVfC6wp9IjJ9u+f+hTA/a7mgo9mNgk++vX
9jCGRiXGowkfLiTf44+uM743hscWFaWgs9/yyjSuT22s5XvW88XsCZlHGDQUUuhV1zP1WxG2A7Qj
U5683Lqltc2IUldy1OOZDdrZrW7mY0Fxl+j+9T5IOo9s7lvCFDYsl9YFl4n2Hc64IIssKqyCYJ0c
BMdH02yvhET24ZmZkeQm4PPKUkOvH6uJb5ZXod7UfRj8wm7Iqb8UlOaUEBmAtleyX4ch5lXJz0aD
zGJqE3up69ngTuk7X4sG+L1jLeTu+ln3siZOURK/rvgl9/qmgqktywx/ErDN2PeLh2/Cx4OkH6zu
P/ZyeaY5WV+g+CMpL0gYYrdMAgrDi5tvxi+GLFvb5vcJsdzzKOLFJIroGUIDnkq/N7xdm3MyPA43
WwJTenICfZFVGw6Jdyo5mCTNPk1pAFCjePE08rmmKz3JX+f1s9jQfffm5a3vvtOsBr+jbf/MlAkS
krATyVLnY9S6IWVg+SjEZp72+msKldAfvjYZ6HGKpC95mz1alEcefM8nxQuo77msZoUr/k3rFSI0
1BEabuoC0WpO7TBeVzu9Ar6ZgjRqDBZD4oUpgAVvnCcUCbfgkBGN1OUzyNH6yK2nz6LRzRddaCfx
Alr6oDs5cwMaCzjaOAxQh/LutAwZhwo+uu+lmKGIxtAWpaw45gxhGmgJ9UtJwqY+tKE3PoqFCfQP
N6TWM0mKx9kbkHnBjuBaexwSaqoQBDnLrF8ZgQjoa6O9uqaHEbxzZJuiG//dKaEXxz1PliU/FkS4
SYaE56sIlDwn06BhKRgin7ZVEwr5IVpMEMQwdOsvvnrploBEl9zmBds7cPMjyqA8WcfgAY9IsmWi
jIXkpcLY3lreDrfzpW8Df/q1nk7u0FvwEy5tUUpK7ud26CiXjY6YucHfWIz+upYMf0gz5VOTGE5E
0rJmtBVehfzPWssToDaccBDx7cRrFPrkKtfAhTp4v596mZfEWXvKbbP8mX2OhC/yyrHtnziHKJWF
D8oTGcsSDYS3VW1uZmaJln7GAAfKWiWu/LqkE6s90gnCINmzNWR69PAnQ6z4VAq9YDhjz0AQXFQ9
iK12+cUqBHwiVH4wafBICDs+Y6QGAJ3aeznqViH9EUWQ19XsMjgVgSjO7uRDHEq5+7whQCaBsGNl
BaYRk8XPRpaY6WtU4ZF3foH7623e/fz8vVqW7k5BNy/C4CYz4klhy6uy/t2CfevQKhXMResOn58V
W3jyW+ayWyKpo25cbIJt21MAXCer94LOo6fhBZlLJmjSmBTWIZlFZ2xMWwFCo1FaKLIw8EH7Oyue
WmCzjU8F2R/NywUUkq14P8890Jy3UrwDR2jmDUNqotGLw8c/dvZ0KO4899t1WeQAWD44nN9IAiT3
ZEtgC04+0cFnagoXgVOR1dzzdS+Ud2piV/yaKtJYnTqjWZhhcrhaKxa+Wl5wL9oX/S2QRSt+D86t
OgiKjdqoSzdwKcLddVH20EEMEhpWet84J9vG5NIzCnH9fjiwSB/auDc0oN9dmiiYkaVB7ZntduGd
IaKF2BfbgJn+HLqtdIy5nAlT+Zzq3CZ0K6vLrWaV0HBqjN+W/ywb9iGZq85HVLTH5lBpc/CfN/c/
UIdredSLoR07HsXFVfwyCAP6MA4Ak2srXa7xEqE3rHJMaSdus11Kawp+lX7IT8Udy7bI2OoShchZ
CZVtgL1Zxd2k5Lq+KfVKG9fdPpiuawgmsyIbyGnfEutxMs3LeQUyVPsaM+DIagkU97yCPuoRBrR4
dacRHbzq2s/P2FE3775M4sMaE2ZwCmfleFNmh0pjGFA3T5aGVfKbG+PnXFKUNNeOaE/hIEgxu66U
MauTcRBeRJ1QOysmXzF28zxR5neHdzNOTzN4K5i/5VSXZwE3vBkh87e4MCXTBr0jq1aidR2BknTs
R1bMfrQRJWkWuj9niBFuskjHEBL1zUmL04/xLDk040AS2r6gCskFdshLmXAW0JLsqW5XvO4EztHE
9xqlOgTT9UrWbFHVzK6LRY99jELwErlGG3DMy2MFZrdtjBPW8IcjA1UAhdFTFrjxDBrWLXOAxQWj
aVXItejWeX0UuCawqkf/rRee+giMt73whkEZNPJcNkEpoKzHW/JafnaagSAvNGYKsnj0jjrAr2Oi
iq2804pdYSve8XNF1i6k9ljiIbswi6Uqn6bxMTIHzSYlh/+9jflCEfRb00RnMsxHaRDxySDf7P70
eApk5kqcSRga9jszQPCJXhNBftwTJ1vNEkYKlfGUk5vQ7H0d6/8rnB1NgKviXZUsXL3ffOan1kc+
Khoo3AHIxEDKbopWFQ2+S0wAd3DNogwWpXi5EgPgAbl1HMCAbM42osfe5jjvZ12i623s6lpgHWfE
r62hW/WMAdSRMDwBbVyAwiAyzaVsZmi4HUvzyTcx8J4BXH6EztSz0B//wfcRP0N1+Uae3B0zesqK
Lmpgi1CJ+5nbff6Hn9juh7wttL5NVisi9byuzs9V4P8qIBo68HHYrmPUy/wkfOXSABngimBAf2pp
hI1Nox2K0c99IP9ZnSYmn26YaaPA2VhSoZKr8sXfv4jMBiLgzLLP/QdEPfXOYSSFYYmyCsX0l6Zc
7Gra8ZVtJkSp6AL6qGuAfDOsIqNJ4n9oiXTZmO7oD3sc1PLWE/yA8fe0pLEvFXxHG1Xz7/Y/o3iF
9YKY+skTvVWKw7AZJzdoZ/VCfPA5gZAYH0EA/tI5DTuX3vGZIgMKxyw+h4c6UA3Oh5md/Dz6mDkQ
M4l654VTStR6I3Wy5sjf7SHU7A+c3zheJ6XBpFrxf6/cmowkZGu7pYD1srU/IwVet79YoWYQt9U6
YucjXZKCc+53gJ4Xp2vOAAWYhEbW+TiXOwjWvtkf3JK4XPxfufFLo6zFYNKAEGtKe4xzUSTE+rn8
uzBHdqFnJCB6Bc0q9npnnbVZr3tpH/L8CBHURsjO4R6Vku102GFj/YhhnapYKNPEqkagl3NZpNs5
gfs3Wgy32a6y+VJDI28WRgU4aQpk0qB4l60ek1mXKE5QBCGXSKFahH3vFgkmd+FKLF0UODxBGHuZ
ZRr3+TUFE9/2jtzU+23xNmL8Xa7A42EFNHTUUEmB18a69ZD39Kx5zbToQZ8/oxFBvpbiPL93fM3Q
9bhA4MBLsALaC0hjn0nK2Yk+7RFxlUMzIiG5W91O+uirtblkogNsivKjYn7KGG44cIs867WGDNaC
Sjc14Zm/K4cMcoyEWx5+vbbMYm4rDloitx+xp44N4RvguyaoWGZpqYbILvUDdFyKgYdssCH2QHaA
lVegbVX6VetuwU7jPwX+gf35iBPtsAQM7QqoMWFGI41Jj5oXeyXnyf1JXCmU6mxasKkNg+KgjgXj
spJJOxolNFYGezmm7lmSXUAqvA/lvQyH2wrFKgcO69v7AkMBOa95NSnP6jwcKlt/kSqOK6Bzql6V
mxETAW6q3AXIiAmpZUT6Xb2dw9l23Z/6THqw7nJ8Z+jan+Z/Y4bNAaEzV8WQdJTtGZLqlCp7awh9
rqC+DPUyhC06xKNbpyJnpinwsuE6q60yrw2zFJZa7zb2XQdjdeIvIAF2yZvkfEy4YJR/oxs7fHci
uf1NS6SgoiScTAFvDbAiFhIpWPCgMgJxMP5TmQBHzlLvsbSwkXPXNll9zJ6stbse7S3Gz9UOQLV2
ABD+hqsKi/IhQXz32GnjXP8iLCz8bGNYxYlWL79XqFb8KDPGXSxIuu3D4As6a7OLbmDnonuUiteK
xKl/NhSxA44R55fm3v25WSJHqs1WSWBMQMec/qP/hfhqZId6VUlg1Z6f5enpt6o0EFtqWd3auPco
Fc7PHeRG+0LbccZHAevdE3kcCaBH/sK1MBqDEBBPlIYoBZK8FLdeIl+SuDscJjWks9IanVW/iEi+
/LoyBCDtJ1kb9pnzxvJ7EW8Onjl7etzwIkUKSsbLkrAh+0HOH6yh2uwvk8+N/hYOgdYycCARWnrB
x8EUtWr1q+QEmeB5wr9WSIl/ytT0kHva/mk2aJBjln7fvTJfjr/nFLYW428XUttVFDlMoL8FYMIV
2ntq3YNxL/j2aYzuS9lBoejmKh0DOrD7WP46jlFy8LrwhWOY/rbafnXdY17/ak0/2OIAjWeCkJJn
Fh8kmljTX6DWrcN6u1b6iNGQEDGbqpdxwl8foe6zxMLcBjtjru7cx3rjhBdwtMFFBYq2TyYLcv87
lM2aQyhTY5ooJMx+2V73VdmhLhBrHQTyB16pFBpb3OgzfKNJ2l0BCgPkEalu+YecdrUh763tnTjp
K+m4lOC7ZIyERu3nnTc6Lq7t10bCeumDuwjDeAU6shAXtoH6q8MYXpKuXTYjOg9MnkuSF7QgIY5v
YcjeuU4EWhVQTM0gORLqB+QzTv50Uie4p0f/lplo6uEeph1PXf8pCnXgVx6y3HFd8VN2cfLGvp8K
TFjV0HCUYBoGqr0L4qi7b3dvA1mHxMD00kRpG+k2BHD5SrtL18OVm2xeArMoNJHRVNChpwnletdJ
9qRYUk8TZnwZ2lV6zG21SwHsd7Sz6Rsyf78jClYhD3fvCYlotQHCdMTSXWQfVHDW1MrxjOIkbazx
lnD6gvniIHF6vTGAx1F8QB+wp+Bw9N8nwSqlCdIuaZQ5mUlRt6UZVW7ScO+bKZEGbqJ83gfB7g33
N2mLhhwJA9O22U0QtjXRieqBmiDhrfLhozWluOcKyl/RZHibJfj9WwELTNXMSo0LdQ1RE3nE37L9
6xtcckNdD/F3W63X8qg5/W0/PGvR24Lf/I3lV+1rYiueClLoYSShh+V+iFFsuadw05qXswTBqm/n
TOtqI+OOgirIh7rGrusyCxGFpx4fxOArCcXmVf/Zk+VkglScS6TWld8CtoFIGC2QhSZ1j/9m1bTV
MyTY4WX7eXEYjHtkt/4xI2aylzJxxhuhGgxMwsqO6z0E1kFT84MTLMDY0CfIAPmNgBeAgo0C8QVa
Xbr7w9pVviM3v6YxeRqyTMk1BSEFRVw20wWHFqJIsatmfzood+M16rmpDtfuqfnOEOsCcGVn4wQk
21BnpBKENIFGGOz+M4/xLNn2K9qdkrLX4RSeohpaIb97TdjtTPiCE2T6KzaeaM2VTOv4nfHubc2E
nz3Y/sp5TDHBzue6NUf+IB3vgSgZYSAIJ8oBU+ijouaSX2eFuLNJQj2O4zz/sBHL6A5DXLEzE3dn
1UkGiKsOdHm7JOokknXL/fM7XgkMLUx+XUAlUeBhOf2clLxShIdSfUJTnOsFsvIWQn3vk21pLifg
HhqfHQtfrqCSj1BgONy9gftfv+6uT2izzBg/k/KtHlj2C41KL5uwMWhuv4X7kvAJniurfjvnEORz
hTvMkVr54Ay+TT+Qvi/h0V4g+K2SmtXDcNU8wq2MWGvauFo1/+KOxF48wZaclqrHYAPOUwnW5t8S
SiXnwn4N04whj6UTLIm3cMOmD/kWqAVkWU05vSrS6RzXCVH6jaD4Ru2hswpe5CXkR3qmf7xRVyoL
5dgLSGZ7JQekHEVuAT0lmTmqVs1sx7nWf840ouSQuywcInwFGuR9rEeZqAZ/vJf0cXVfRfSiWIl1
co/mK2U3w8Kx6FGyE5komfQ/eWpJSkLM0TqTNBE2kH8gmsp07wWGqQj6gh4XjCI9lKmlTgwpJ8GZ
TiK+TcHdqSPQ6nP/9YkpsnO7bRaA8CnwhFRCNZQWQHsYMObqdIDslxQwbLGv9+/ZJBrngdPOjVdn
eAZtEOBIevAJqEFoWmSDr/ET3AKeJm3FaFrsr+qmMVLpUnBFQprFgeOBfKr5u7IW4lZHFS8LsQP4
19TC0Bo8rdoeSJCUbtdqb47YbU3pKSFPlUWYLo/QOiPjZvaXlK3B6XdA8iU62gIf8qZ1Z36lRDxA
M3cH4ClM7dh/Oh0z48C+gP6Y929wkWU2LRAVX+K84KZSYbVURDjddO7ZROTdZS8TIim02YaCj7ck
sUy9rD7+VUrZbMEjrzVjUHxfw++JOMVKzoV6u5aG7G+i/IkKTngedRebRJKWR6pnou6BQuDk7sRk
JL6GQBiTULjmTtstl9jMSZODl/Ck1TQwTj1jLmsD6cIfw70xKovrCOnEYaBlFGGTbWlAfmEsx48l
t2WhkcyzZTAWYLF6hplbVBl32RiEledMi2F+b+PcJAjOobBxiN/7AMt0flIGjjn05CCF2zv/B0/7
34K/LvRMT4LmqJkzuEP/0m2WhgF4CfcuGFImd4N1MlGW+vA251WRwqs8AUSkIXFhyMMyLPP4SX81
ahyItQqIU1xrstxqNDZjNVMJeo6DQ4oI29QDClhKnBT3dLDb22V5poN0T2hE9oHEEpBOnTBdUqqR
zl3QD/nhC9IgVu2Ctd4QYVIsK63qMu1WGDOGBA0O8rp8dQ2U788FkraRh0Gp8WcrBN/DBKzvupkF
LB+5RkDES0oDdKoP8lnX5veXweN8KT4DOVloAi61xySRu0EQAo9xYUOp/2vjYGL87NsMEFbRRilO
qpsiO2jPqdE9xVg1pv7g2NB8JJI9dmfDdsTi1K8pdXAPg6z8hBtccP2QkIXOWBEuHB9HxCabBQT4
cHH/7vrrZsKiJT4f+1A3pNv++vJ9Q0BkcOlizp4lJICPGzqlU6brpvm20ib7ZeO19vS2HzlgRv7s
8P8sT7ZKx3EtZarhA/crzYMCoeHzH3mvosNS1wN/x8TIjjAA6tbG89pByjhkkfCOSN7gwq5e3Ard
XkvdwKy3hRqDm3Im8I+NrF8HuAcpKSvjSRX0uur18IMWWBGIggeXwPbAF8+SkQOS6gVxUIpX/6bP
JGxFUxqMQA4M/S5Q63zRhJr9XOLTCLjZBriy/q293/XSb92HMcrh16APFAn3dPr8aRFSN91nQ3Bv
XP0JKHB+Q3IFauzJSamiFTso7KlXm82KXdy6PHgFELHwFIXwlfqnN3E4XH6oOlOQoHOs8Ry0Hush
DLmQF0HRNIHm+/crFfbjLgqlgmWKDx26dXPs5nyvNzgRfioQFpDNrX975fnYKpC1h/hFNtH8SFo4
2pLZXE4OATcdci6s5KC7IrbFotdsEs2LRdRMq0/3Q2MlAXH2Bum8m7uefvAL9DbPydli6bDvvlXc
/eLWeId9V7UqNJvt/Nb2QhEb3flknljPJaQ1zRz3a53v7UIl4ThmNOnDdC+7vJeuNEutrn3oqK5C
l9y4prXTDeDg4f6/LYTMbh8jCq25bCVp9C/2FU66dDnECq7i4mxheZEFgcpaFRT/K0zq+J19Qa8Q
DCvWad76C6+c75lYkFcHQQC8G6jjnnCRSIv9Mm1WfQfFma43AkCXzWcVkk4BlLnFnsNdF7V+lvJN
ugTRPWlE/MKi24DnS8EtPcw+ljBdNlC7RtNW9/sIr/pEk4v0Za29B5fVIx/29H4P1IAS2ntECEWd
S6JoifMFMO7f+mf/w/VwX/EYt4JgmYwcy63DP8v/R9ZgvD9FsVXevi+pS3fjUlMRm+G3r0QahOG+
f5oEokViZz50Z+F2QWefQcBTi7fIA27Yd6c/Za5PujqeGyiYvdxg7bJdC1d3dPwpnVRS61vORZ2m
lgMkGOTkuctrAn9ZUyktVipz2swwZzmk6bBo142JbHwQSghb/Q2Tzee1+Jjd5E8whtA7I99JqFTx
sikCCBzQwcx8ZQwe5mSI5+WFPphC2JxxErDvF7tyHMDOTVVwNdFqvRy1TCH4UZfTa6ggepUQgF7B
3DHbjdGvoJ1Smeava7/y51xpD1rG0bp9tXKL4rgfQlpJKyP26PVPcbgv3wo9uD9uKVQsmVm5E748
MJgUVSJLa0NB5fH9oQystyaRBX62IRimnuzt9ddWSB5GNQewr5cf67GCiDXTMky/lKldQPlmNWEi
sLLIn6BWdCjzWR0t3yPshwKPhBHMIEBGLp0+Qds8UznW06BkMVEuZhXSGSNgrrfMTIrnL4kqkcyZ
iEdriwcWd4fSZk5CUiIUuoJOeuVljQsq+uerg/zWuotojM+EylWN4jE5a9Z6dAQ9fyFDUJToWSGu
yvmI+xpzX85yDE6Gtr/0W/3eVpmZ9vk2VKV9xLc+Lbn2SKIypjhcGqanvBZ1HnZKKM8eSAXpTcYh
FZpfpGatZpufkvRaogwaJpkpBh9Cw8wHiruQqaefEUiN7QocAQ5+WTICA33e3fLPKGfxHchvxCI3
KeMLzv6qTE0F+OuxDJva3041v1dWrNeiuS6bMS8khf+5qzQUCD3pCyT/XRhVGDqlKbRzTl1BQTfP
L8OVCmtih1NDe+Dm//Gc7fJ6exGlbZotD48ZEx/5YeMuxfV656eTSiPD9a+bsX5sF2VUEjHKhI7I
x5l7ilgNHwWYHUghay01msEAic0rHmxougqNzZMP+EyM6884o9PDLF7/Her/ny15IUYkwLcIrFeT
PARau/A/Ue6gtKf4zeIDDAaytRQG8Vy4UOwkFFH4pkeXLeJjWBdf1WS5kOltzVo1omKLMyWd4Zpb
G6fpEA64/8DxFeNb9SeWL+lq9GqHv9gB0d7X7BuZgcya84kFqyV9T+joqyu2XxO9ZBsY6qAL1kx0
MOWwGjVo/DptkN1p6nCBfDa+Qu7T2j6rEM2F/fyyH2ohXjBOgrjaHsMSJUB3nOC2S5YPfap2CoPP
p6C4aU98pg4O6ZxerkTX/LawuHYVJLwB7N38IYCLoCbYJBtNlxwFcpI75XnFFKE6MOtIVoIRDiK5
pGq/9IZlXhE5jD1tSSbWI+MCY7cvRogfxTjYwq4F88mMfEuMbTl/a9FJm+3AMZmhx2TqI+VrGmoQ
PLXJ24F37uPy/m1wEzdT2DQqbahWLUaTw5a6aRj/Yp/zc/SGQiLCUOaWTN3bnjN/ofFYfRkNZf36
aw8s48AIdZ+LhL/Ff0RsVpDQ0WbZaIZmGE8K03gV039pUa5e5+YXeYE3I4y7iI8b7UQh7SrdESlk
VO0MsFVNIcVSscGYFpNL052KcuyN+sbVMMBmRAajvzWMOPZLexMlXhZCX1mINCTlizV30SHJkBfh
IUfCZeK/75UNXV4iunHvTgxHXjn2RtbV6TgQoN6U3WBfGLS1AvQBsOtX6UtLlxjRsGpgOkPB9aqI
rBUtfyedpAD8z4xp3v3gU9Ju016bdIy5d5G3Qv9htaE0YKeRpPZsEUBHr8edkkOR5d1za/0Xt628
IeMVmIdusm+etpdpc0kmTjR2tciP8SftsMiW/lEPB6TwER7B/2A03tbfHan9qBENWf0Y5vLVMa/d
3WhRPbRclGn8a2rkoSKF+5j0+2l+4ZPN7dhiGkPnAtkSwbJStVVnvFJCXW76ifAIBC+e0faJ+idh
j4BSRIfpXuKWeNmJBk9iqbVMhEGqyC9uBSGKoDFb1CT5xDCtjAlzJ+ENpj3vdUIDi0REI3+aJvAX
mX/rsziCXoCEiUuf9MmBvL7Hk3v4UkoQHWPtd3kvJvUGevOj9gyTwB9C8q2DC37zL17t28Z+a107
6fT4NPvnQZpnB451bQupIdeLgXZ8sdy1pFzkBdOUuCaN1EQiDCAa+StTYUHiE9LhPKrweXzvvhvZ
YZ0e7QJTS9KjxuCN7SSqbpatoRLKMsMIcpL+y29v0e7lMq4DMamshQrxiluoquDNP4rnH3BNJW63
gVEEAPvhRBoS2CtZjxJxvV7N40mdtGL93POFQosVKagdhe0YHQ9uRdrr+P2DRq8/0BBeXqqS4PS1
hFKAtFonaZrqMJzq4TU/IcJiPeRS76+ljGKRE4lwa9MdwvDdb0v1sLmlGXyGlG6leWXV5tGdvxfy
WCquKH7WFG0QBcfFmOoXgG+RElIF/PMJSaH5CDpmJR9mlCcSb6BZvXC1du1KazF7W774ke7krwPk
38cDApU3gxYFAQioFBV/SGiadVQoBsS3vlRFvnTQeviJd9iJnwMDADulXkZJs8HY2GYWtvxEGHVP
kyFSp3r2LXeOhn8KtgCvAlnhbRoYraHvued3Lf0cNzI5vV9m54im+AvJl1x/b7konyioPYzhr33L
H2GsDQctoskLZji4oCuBgCYoZNmdtmq7z21qYuKqXBQzL4wvcclm/LdnnDEhSj5KrF9BqB3wLV27
yYIW/AlTjSXPxFYcglUekCCsZDGXOE4eYVzgSuYdR+YwEJFLemQ7cJE11c9UPXdFnj88NEQ5KLwk
G/1nqOeKyOeHV+5Ho1ChbaGx83X+CubXESESHjqk471KKAleFQwOEWJv3W7cXV7TPGxzIGwUboRO
E7aKkcrmguMRgWm4flntV/02gTmmuXhbzZiTe+5njOmeGleeenw/Qd2ncMoRuPlfutzr9vp4r7bc
4umhQ/+u5qhLVzBl2t8mowAlAmVWhKzmKQZHWRjwFQx/BXG88yeUw1QxESS33l8Sol7nKBU217N6
c2mkIW+iofmfcu4cCwIhNvt9eSb+I/knWLfEF5wzfYEwZfu30eUaV9TQY0PQ9cVSvsA/SH0UEjly
o/MhhaO3EtTljf/oaPRFOHTlCvJtz914KdbAO2llwFJATiiupWAZ5cxy0pcW+q+XNVdLE1Ndt93T
VtRutgkAf4om2b8DXmTwhaB3OJxxk+ap6vDcOPiEYEV3KHNMZgR2nykNSoHktxLXo9A3yaDtWR+8
z4yhjYDCUPBVXoREF9xLuWjzzdRQUFuhAJKGIk5117fL4KhZV2TJHUwBnSgP++gSGPOKCCVAE5Km
AjQUQL/xSOo3v7lCKBKdMxrDSyoqwTD6OCLcO30KXSYHBER+t7cU28pkQqifuJ1kGIlPwGt6T7Q4
+v/xUWdnlCXiSiq9SMdj9sWt4lkp6yCvrBC0tXS/IZZ6GrndMZqdQPktm/e29eLmeze4ky6rDvOs
xXlQ8LU0qDULbKdmqReX8oszdgsmownJd7x0TFkxp41joV9aPkhYpEBjqo9aIwGFGO49kV8xjfTH
BIYfsuMN++HAZ45K4CMAH3mHfkdVUzoj/wPQ1KkGco4AB82hl4Zd7477NzbyIkbMgxPOBDQk/+bC
ZeJLM20B/sBOjAeQ1Lzu59VOnmmHJpKEhgAwCDy/BbB+mWbfch+HaDRgynLOc1A23J00RA6aFpDt
cTbmelGQL6do/dD5JzUIABj5YG0q315ihcDY9xfOKhlEaSw7qSZEspl5GC6xgQuWODRl6htbct3O
wjcz2MQdr+YZO/5OpYvL1b0vlNSP5XfAxdPVHSTzHbs8e0wQv1Bj4e5Mbyn1camH8Pc0DeIgQK63
vBPRFcBbwZ8eIANRKgTIXGgUd1RBpX3d+qYEUdk1VEwWnbKCL0j6Yi/chnsXG+EhphVZ55tYpCln
bRSSjHE80+xIK79IpDZtT7yjCA1oQRsgpEH6D/KiCBuMeXRCYpPB+QPx8LciRKOPoM0cKux2O807
J4+CjPdbNbj6DYS7LVN8eaOveR5Cl+PSASpqWbw+rArFXAVYM3OqExTwduU80XIQ3ZJiIDGqXgVx
dRenkbarFGPuEmBJJsocARxyT1OmqGVpkDEi7YrZ4F2+RbzdSH18aajobmmijWtO6w8OjaX3fTnH
Gu9RvZ3t94/kv7p+kmvvg4YFkuO1eMbF8VhdN/2NpJCVY7wl7spxTCksfuukGDAgxM65vEahvKRJ
1RPENHeEHZEAMQO8U5kL2uj74qMmwqqKeBX0k14b1kADq7r2r6grUjlFjBxxhlq/uzOLt3/XjN2d
vC+EC++NVYMS2JH1mQjfBd3UEacAsxdEoglgDgvi6gt0catcng4E6YUifaA2/q4bUHKxJPbTZBEl
DjXFIBXt8WKVzKMX9/QDY4W7+Y+zMVM21oGc/sJWaGOBWUjX7c+dpqF61CXFovvddSvkuV5baEhn
5wmfhF9nKaQX1wUTap2NGLYQPT/FbrR6GksFnifdYqh3ff6OoTE1i9bUB74RPE76qEeb48sjbt72
loChHd13NJAqlGnxtiDVolpqO7tC/wCDvjkWSsNiHCW2LXhLqZpqyfUctMvh8vMdBNhzfZYClI8I
cMFk6qIRclW1zQq+VMLbIz27ly/je1bObBAEvNsCS5lnT87Nn9A8jRzBXs3Nw5XI7i9nW3ZO3ubJ
WO/B8IHC55B3VOyH9hSAKgRYEXlP8MCDcUhFZcjM4/XMWbcYKF0nnDfRQzr0VlzYISFW846UhIFt
tgJfb2n/mrNKl/tBz96sRvURqfujdTUiHn3mHhGJmtgCs6Tl5OwVKQ5mCUXJXgpq5gXFHY2CqWUx
KWWNwZ4sYjICTp2EgJutJDmbPkt7EvykpbkhzkP3GlCJ054yaZOahhIA3KW2g77se1AvFFnecklE
rudqNodiDmAiDfwIeomchadYx0ZERqN5JZRLG7757hQxYeZceIvynX+P2462/KiHET1ainp4ii1L
zh714COO0LR0p92eUIWGDJrbQdJZmekH5kE5FWvGOD2UhfqIVwgsWGC2mxzbDJSuLo42BwqNcwsV
bhPJ9jh8jdiWZwR9Qk9Uyt4VuymisPe/7u+D0jFsIxDn0veeLrmQP/e5hEOX1yrEMoD85onvYqA3
+AnsMNVZljGUlTrc87wcukiwKiioIcsEF9EJLaEFBRghCY1MCpRAUFsX4boliCP6zmMA8ra8Yv0a
if2LvHXon+Nhm4SlERMP3JkgeCHTvReEMsFRcWhZ0f2r7AiNhRdZnM6wUsE7jS4f5WFm5WML23hv
asPVERzELjUMTDV3Bs2+YTDXyYh7OIZlyFHnxp0IlQPUu8TLDrKdniRHnauUKDw481ql9nMnEDsS
13TdRjmAOFQTseTwXQ7bys9ygM7OKlHfDzmJi2wKoAoJXl5Yr5d8aoGrSluz5++H1q4kNYpprH+Z
0/YwtHeaO2Uira6NX6lgX07e7BiVvaiITaNyjbem43n11Lkbxcf6q6318rOgj9R1+qjFwbsL4uLr
9zclO1RbdKfUbaOiNq6ayHNIMN739Sj8Z+WdMrxYxUKnuqn1q4c3kW90aqFaC4A9jsToAGHR3Z+/
zCcNpX3zEAzqEUPyFy5ZWigzDr9mnenf65KVFmqm74LWnG2BiTgY46AeC799xKbpgWgY556G4jUi
jz0fd8zGVTvRjVwbKC6vavDAxQEvXtK2RatPWJubHaXDYAQHi0DR8/BW1j355sRcqStwo/4LkAfA
QNARJN7bNe6SlZiTqy4xn4goO46iWjakR1n1ODaX2W9rpsVrvJn+9qGeZX4Ozv82EGeHdNXunQgA
gUAhimmUS97PBKBYHw8cszafWAltyY5rWlkM+Ens/2uluCklMTys1gyhOtTZFc2Cs/vYr/eUP2Ua
x3WuawwbdWsrX+078mGK4SSm0rUsZL8WK5zDjOgkNzQ1LdBut0ElWg3oZLI1IC89l+bCwYaun39x
LtPYQMqGtBlEWqctpLZ9j1aM2ubSHhzvJoxvBhnPAM6b9mEOxMtF2BNn0zwCw2EFDzcgmvPOqPvu
vAlx3xtQbQCrKGi4pwcRQH32bXcbhbCKiABmXAU1P5SCq/ZoRGbV+xV+Z8M+cV/1YO9xtKYP8hTv
94RBKiIWer4oJ/ZcEQaZtoICLDeHbPFp2hqSVafpeP0oNLe+b28zwcULQGetdmapN5CSFT2gtuU1
coVtoYsk66BOPqoFDy4j/eYoStcmBMkVisVKAqz3Tl+KXy1ozoTekcSBoMXVvwTkD37VQpWcdSXo
UXk9Vo6mM2YO20BvnsmCFqb+QfwKx0OdQ3HRPKcRa/5r4Hc7l7evnjN/7vIE3RpO67HquV7jmCkh
AF6dtwKhii1Dr49uwp23l+xmD0lsHpkCFLHJd00XSjR1CBYC6QnN+23LoV1NsdHxCGHu0aj9wFVV
3qWLuf8mpGXmWnlnHO3Yqq15O9cvapgr2DG/AZ3DQTeSibPIaKf05WuRqnMPX95i3OBoxw0MUAxR
t7HIQuswpL7R6AFZsbDbyZRNZhoDYYfVUlv7GAnAgaOvsNa0X9vnI52bTtYVI3BDNim9e6DdvsKt
8FM0ektPTuYvfWxmT6vmkdfyPUHXeXMlS/jWywsY7moY3SlpOaEiwF4Z8smox46GoesTdvBOhddv
WGGv5hOoa+xq3zC26jppVLf/hl1oo4h0YjsOC7SMY9rTndynohn9zwCb+FNCCKqmrc05+x3jGBGc
jLYi/Gv7yygHS7nFRWSqAN1Ss6GLbrT6ZCpdnxSwUvFZPa7CHG5L9yOJonlCVT7udhyK/zlRqiob
92kXTGZ/uj2m41kLVHPW99DDaPl6A92PJbT892+kQmjoDiBRAFyvNFs51o1tPx3kIwMaNJ1cE0+N
QSF2DwMegJlKzAYODBwVsiegMf8cRx5MioNlS7e+CUf5zNZT9vjihKc3qJCxJEYpw3z7tYoefeUs
YWlaZh82nlvGvB497GOb9wgLLEnRlsYyWNY9zl1hGmsTE/39WRybDk6e8oBlEZzUD4ItRMGGM7iL
GbbAXUQeMokAfPc+JAY/o/BXemCrgxB8yCcqxT9A3zP3j5IJUnAJG/FbKrKZV3CEd3r9WbQgIENr
QlgRDIh6R+6YeWiHsN8N2NZJPEf/gEs31iD7GXUGiCPFt88bruzBzp5KpGCiyPnMDs1ZildT276+
audkUCpCubQNqZx9C1Bpe6LyVWdxAKzJRfCLB7V8Vqcx9IHIHPTiiXPZ78WCOVGhUvxksvq7Dpk/
u46zsItgQ1U6O55BIYV+zLf/m/WkvDprn50S3YaOGFKp81c8TC9MaH1t9kT2x/g1xOQXZOIU3QgV
eSTrCDk1lfz4MmbvCzCxyV5hbu9Dtj9ReV5Tpl+y9SF5acAbqpbL8lfSftpISy+dFPT8mzse1BRe
xf96JWTUkz1p0vapLhmSa4rc833CrDn+ifwzjdM+ivTEAZaX/OuwaGe3pklZ0DOyUjVRs0hxN5rU
frxn62fAV8giwgN1G1DmyqFzaEjUASZOGV3eEeA7Ruxema/PxSH10xUYgOQaTqN/N2Vj9doMNvoW
2o2HqGFnaL34QfjP/zwi8aVtW9ONT8q9vZXYERV4bFR4n0dWo5oeATA2xDW81lhJ0ipD3MoVEwPl
jB+RaZGPqcQ7Vf3SsS8JosCLsIG6AmXXleds97sWUybbrPcTWcZjYVkVr+0ruiYcz6lGHsWHENOe
jnVlmar+FG6eFDzllNSEDxPWo+pMsxxbB6jyZ8KOnXxivDFwQq0QtYMI01vEyvoZcfF6HqaCuunc
tFLnhZEmVPI1xFgCBOO0cAHaFavrksDRHYqiIASBl7qZRDdaYdJ7T+uTi3UKDn7Z5F6/gtBgAxl2
CUPla0T0Dr4p5762m+gAM30smLjhDuWpXmYKdMfPxBmw8XEk4+1hDG/wR39+W02JkQU2lzd0OOqS
BGLUlqxW7yjYF4A06PBL7edYWQ7JcrSJ98lBa7MAUxj5uYeUS1EVaGjlHFBOEzrXeg7sivd4qA3X
62kmtpFIfKFdIxFRNvSceiKJeT0z4aFHcVxsQ77IPDp4aJsdbaukNK+4AZkd2PbYjtJcvqqRTe2+
yv3Vj8QppSklgqpjiahi9ed9+NocW7tf06XupMVJMQZdgm5S5K46X8t0YEZiPryOxz5LoOOActC9
b1grzWlsI0lVXITHIO8wWSoisOTIOHSwbpfeQ35a0ui2H85UQOazdftyRND7DOgfBJ1Unrvnl8SB
WhdziaUygmMA5p8jcHL91MoJ+X46fwbPVt1GrNRkkAUSHUTfmS+D5HtEDbTFNOU6oByZlZOcXPxa
OnHLCYXnYwhZ71FCfXwQLDFbnH/omSQBhl9EBR2DSFvMRV5gmh9wPae3opmoctnhrLXr2MZRZ6/m
Jqi7wZBIkeQn7c6V536bWEW+vogxZ9i8HBNppEZHK73oPek0akfKEjjOHw42uBbviMKDFYhnGHs3
MtvLF2wzH8olEbttAgd9dCE0YevthiCELGLcj0yhbNi+naaMypxRxbuHqra1Ez4RzIodSyZsF87u
yn5XXRNruEiwFB52gCk4oNlVsqT5yawbMXp2RnBpYZAgAG61YGoxcQ984ve1GU371/4W3m4Wxhsz
7tI6ljwqmG85jCw6/GdYGyy32e56gJXseibB/bZ7QUj7QkxKtiynPJffdB/p2srPEjl/+bPQl2AK
O6y4LEQ4vDHMkjmRiZn/YC6EMgZo1e1zM2lG3M+JDnBDlzYIptTji9h2n8ntsltdUgNrMV5FMWi+
B5931biYWo3cV0XopPpa7AzpBY1DWrLXdY0HD9ZJ58WetT2abltb43xc5ZSDTe5Cgyg1zsvHSkYy
wR7ncQza9y69AsinP6cAzRvq3fgnf+ZRNZYplRNBK6suOcOYzlvW02idUd49JMwby04CTBjI71ni
CCVRF3Y1H/xWKJbXrAFhYq9ucIZehMG48NR8VO0OPfhvWAJLrNGZObJZpueDSIWs4s0Y4FRchY2D
cyLqVOeCH4OGbooWlco/yd/CfAu5gjr1PEc5GGy3X+0IVL+mIn5v9gyTsRw7YQklLHcHstvs7KjD
DO2pnz+yPz0rSbaI0ENSeEGX/aagIe6lqqjRco+j9412VG+u+GpxJB2vbj0Kx8nXXCLrSy/i/Kwa
430rIclKJUFORAhYZudCAPDZxbYy9jT+T5cPm/qraNxQ3GPJSp8Tbr51VqQiK2/5ABrak+r4jCzZ
ezmiGEZZqEtOs8xnURRaXHTQyFIx4vPKjwzmg6V31qd7R5j3J5UPU9VKVIRL1Cqg+nq7FCfNTmPK
ikRvlaNzxqzT0iAwRhshe1CyvW7cZE/pxWKYO7NpFL8Y+XIo4chaZClpHd1+mG+YUFeVebORtU2C
cKBTLbIVmM88W1TjzmKorvZD42WJGVyNF8hN5Cuom2IYnrkQ8jT7IztBUdhiQyZrn4g1IWOViXNX
36wHyla/aM31fYmgGN5ZMT3roRz/8Dflh6hBVmPsBCzomJUdOW2tkVpNGhQAQw6ZSsq3rpkSxayE
/CF2Ddmmo1lJx0TWef6ypjy5QRMs45yAl61DsBwov05P/pCO4SnnmqvKNMUxzX+pqEnDV6gsToRE
/EPWoybiqed2R0tW6WhVyCjkm7eSuf4cbRS9CukRGrMZyk7AJJgUoH9QLcXV53f3iJkkQvErg+7y
bt5g+qv3nhNGFinfIhKEm8DD4Qq6CEqHNhYizRnlpNBKKriUiqkseG/lFzT8Xb5GP1RR2RKkBa0H
O2H1po6yKft6sGrFDUo2SuYEN0COiyJKODnBi2Fu/L7xFGgLCHsGBpmmRO6hkC2OEXh/RRiYq6SY
c3alcZesq5H/Ed9my3iYaNMwlgzxmCwhK6IU0P5KeDNXBs/G4Y8FM+WnbxgW1pq9Opvt/EFCMwzf
o4YAT/mncpLMOHhBolF5yBcZzx5+qNBv5JjP2cFD2zeX8OPNx56RlxGTmB6C0dBGdWWJEnxxnsWD
Zuc0Sgj5p6MygYh/hoS4vzBJFCjRImN4Eb6gy8ylToZ92fkLz2Fog88Zt45yWIPsBkGdgj98wLgb
15J9eTCzPn+v1zGXp09A/fx/3EyNWaOZEgQcJL8Eh2iYo1aBEDaMcrCWhNYYLSSi0mKDSlqOyCD6
qfPOOtJZEnjcyWknzpsVF41rZEv5runeE6HH565iqIx3cIPVZPGsxoyZ4uEdOAx4htT+MPpo1GCt
9ipMV+YZi7Ubxf7yywP4f4XRZcbXwFOuSxnOuShRJbaVy3DNg6phanw066/1PwbrUk4uTXz+Bmqv
Q6d4AfrFne2c4qSB7cLO9BVTLXu+yB7zoDrGDlm7hS3lZlToLEfUoFznqZ3tZA1JPCsmI+FfhExq
M8oU3LPh+n6413G4D6U3/g9G98IvpQ29l1LwG0e1mYLNqg5r6fchhMJ7LLTJQ+hswi8KceEJKz7a
V+Q6vFIqvc8uUzk6x4qMAQJlClOy/1BUMT6+Hms9Dd9ZqfvoJThxPpOhQ1CjWvUKexX8Hp6hofSY
SbewLIJGPFNxSp3lF5P73SSTQRVlbBRWz1mShf2gbWYNIe0CxAgV4ZEtyl2AgMLrKNDxfpenpJED
kn/o9MFy6t9HruSE6xP374lxsb07w42wjOBxQ0oWCaiFzin1KrSp65Rb+ZRv1jBTFwC03KhEX2mw
QcWZz3Nsv+jYNXLZPPeEV8m/GCMuzpxW/oBhZ7+I/tAmiHLpIffkh8W6e83IT/7AqMvHla2KkxXS
YpfkW6M2ATMD/Dq9/VfCuEhlRPX7h1v21v/o/DYShEoekvOr9ZKd0dBmDcJ3a0mLJzVAa3KV+Yfj
hbPsyjjLVZU3IjmfL62/f2seSDqJo96AaUWJw4I+KEVrm4CjeXWwewROrK1tkM8kNXXiYXu51tCX
kGLuqAHGTlXDy6dfe/Gv82vp53UfNbV6iUxoP9bObxpgtaC+tGB2BQVD2d/SRGSg1UlBkraFmh2K
W9nq8DDAC0Ct34+9mWiq/F7N6xkIf+Y4Tfr9jMBRaXibBqNvpBGmttXn0tJYLydk2A+F5npeuaZk
CIfnWfAJgu70ZdkzIzmSU+4uCpAOlXZqhDGRW/vbLJ+3H19PZp8b/PUxWmYjui5Bb0gqfgy4kXjs
dQxvdEjFNKqnoxsDlxkpXTP2jIBvrUVESMbuRu6TnhTUgrj754M0XETuBviG8KEQj7o9vaEg4ioH
wNpx0YOJiIUqbCae+zzQpPqv2sm1o6WpepvmVWQlO4H7+hmURucyycnWdRYNxtVrQybOshDhS2tV
1VnOOLvlr9OpNXhmMgOOwixmL63D5vIiJpEqQZyYZyloXJ7lQVusq+Y/WBHsWYiwZ3yJ6jFFw62k
dTVSkiPXl4qAK4sbn3pPBPLJXruLdSDhldly8FGS7zBw8TZSj6TCAYDamKs4QR3OXwpEHZGZhjm3
3bw2x87xUUHBTxCxTPjTRbWzcf3zo/hsa5wk2oFBhLeZMPfxKvAnLqr6kWwbMk4IMti0OTvsXQmA
932KNBLrEYVyUfk0u521FZtBrQhlRyxCqufU0wyQet20tAsJ4uG9l7j1kk4u7jxui4NgFBAXx5yU
XjC/2v5KSk4zRHr3sLBGj4L66+sW/6vTMVojV/4aEEnU6joT/01NgCmWfWJ/Hku+00lfwAes/Zkn
JVPbNu2OqhxyCYLdoAiFFTf4CpMGfUh2q/MOQlg0PnFthRJif0izCMM5Blv3I9P0O+3/sDJz6GmC
6MtkCPUgkvkcRQ9Nwd51XBU0Dp9cMNrvsywDDcMo3leLISPn2Z2nKq4CaV+oqVE2+IjNMu8+s0Ix
Ui29fk58dnv6IebGyD01ievVzRqymwGRR70nB37bYBez75foeOQEDiDELZvwwruSeGQSf1fflaVO
jNkA0D9hy6JNIwnFCKzpqzC3wfh2Zy6aaJaxeMIweC/KRwU/nQeUelXiOQr0jfc/E73dyYWUnDDH
tOvgbOydxb8IR/lc8gQ+yHvzitonMMp51nCsQJHjAj+lqyp4fo4GEraWmL82TMwzbOT3TvrVA0ks
zuQ3FEkT9e5tpCY5P1dwPVlbrl4KXCB9kmqdmA1JcJLM0jM5d44hgtruS4PoTDQ4DF9hkWQ0MwR3
7lWJa20LNmTb8X9/sGta6ky98jcPty2gFkp9EwcIutI8ZwSCNOy9hMrGseY5S/GO+9VQOLDTWJf6
p846KunCAmywTspNroo5fF8ceZbjPR3h8nxJ/Hko83/yuPa2GZCFj42WlC2kB3q90dQNk/tocQpK
Q/8t+HvObwTJ/win7XK+WEGyLoCIdvCGxb7tIGFPy8Yit5F1Et7zn2AVchMHJW17ZbPWAnnrHeo2
8NCTzRb+CBnOigBZOmV0ZzjZ+nvU0Wd1eVhM2wUYwyUtQhUFx7CfQ2gNE/x/75pGM6NTdX7BEAj2
o9hv3w5Cuw7ifn1ppsDlRJHE9g3gB/AxB6h3EvyM03VgEb7D4PEcLjGR9MeRjkSDxFNHDEwWwAQ0
8mq3mC9s7LC9RCLzIWxUTfxIwpcagLppyJdKG5OG/+7z6K+4qtQv5ai14cHRX0LtnTkQ9QnSGQAR
HTRl9b9XXFoEQwPItaOTPHNaGXcN9F8p0PYhqD67cH8ypKr1XZUOfOvwG3V8TSUZ/PZkleX5I1lj
P/0zhCNQ9PGbJH5z1tBQhX9p06tHqTMfQDvNek5VcZazmhSifT5zu8Mw723bO0ED6DmzeLIqo+Mi
BT50vXLWFcwqWhGJQX18H+3bSAL+CPtgxDWhM8XNgPFNEdmSsLPHCaOPKJpEoL3Njb0GP78uNSgr
KsIaNM0TXo6Y3FZppoHaB3it8rG/sGlCi++VGyhBnxtJoyhFbq4te7Y9nqOzzxqnmxIAUGnj7LlN
H5Zp4ggLB6Qnusabgano0KtBDs4tC3hK4reOc5bFQBthjJOORJ3UXUBAFfwE433/5iyqw/v5C+cS
Au4gUjbx7jUFcXFLae98ZllQKAnNLlAJAr3tZphVAasAHZjGQuqVSbOWtbI0+lhWsqMy5btMHkY9
rxDNwkzJTsATnEA7xfLjoWdWj9iyg+LpiekfNfoM2PJasBDpGSDE43BpyKyTPwWJ1TTyGJMwvzyu
dT5ufL+T4RwRJWGqB7uMWXMv+M09LuW1sNsvPZYfj5yXMGrkajgSnMZdcJhWgbXTVkdQtyUmfCLI
muDriPM9wJHcdPfo7qT2VFzSZrc9KayPa5W9Lh9wEAKDztgHMtn+Zbtf0Ibb3LHEhltuiD6P1sjv
IPfn1KYUj+GcNnFV0RhRhkOArpxhjmh9J2MHIN/F9pTPWltA+2ykYOjt/hBQ/MEhaaO5huRf5tF+
AWAlcULOvykMkcFRvZS8O28G++FjMkbp/ugZR36QIHWhiUhLv445GF22kIBvyuHgizVydFG197/T
IekNQe7Uw1E8CLooGwqBBrhsyT25GSz/Krvxsj+IZfHGg8aCjFOXaTKdmxtTNWCbOLlgrkJ64DQk
BoXpubtBhPVZzFZWaaWj+n2lHd5ZcsgFbrY8obnr2Hc+LOiHGgRj4t+xxa6zSdmzEnycIMYzBtWS
4nQrDVz5SZEEFEUT07UHt53qoly0Moydj5ncFhlaeR2+vhlkHHUk9yqR0vycoE49Sq28qEYeO8Lt
XTgho3JQ38IkT8rt4GUtgTAe5PqLO7JgpOmiVF51J7PnUybPIoYyYhyF6a/6mitgAlfO+jg+eXPI
2GPT+0iShaBz6DpDEt+ZxSB2MZVwCaHyPbwEIx+oIrzFUjaAeodkqUkUFP4VEUt2QMTzT4szpNqu
I5p6jU901KsvU08POXt7x/HJfvwr+A1R2Qcd+1pAgnNa7cIFPSOCAfYx0yHgFfFKVqMS1MuwrFGS
CvJFBHO7tvD20bTkCPc54aKRKet5d1HWywsELH4BCoCivTxzFpT+ML5I2zi6Z9IseMddtsMoDUqB
8reBBC90FAiIuDqn2/SfPYO2dCbl3Im+TeqKarQLmRKF3+iGjbxUJrnL8DdpLIcPsG6CUHLFKKp0
S0+2PFVI8Po16E4EX+My/A3VmBYeBxPBS8aw4T7UiVV9l1FoZa9+TjbQuuCd+q6yTQ/ZZ2ScRefl
pKbq/NtsmRPH8EPN6wvv4P614DNGDvOJCMyT4dR0OJjItl0ZtKMCNk1fieuo5QZ1zHxScSeUF1jn
BRu9s5UxvhgzL3bwF7EZlg70Fh1bFD0TY+HiUogmfsqo7AeR+zYKgqVRuuAVFsG/SC8690w6t0P/
MZgcWPzdBMvkZEQamjJQxBVmm6Fv9XPKcXQrLt8IwJ+udfsuXapWQEFtUtDI6PLGFawMYmGYbE8t
Nkiz4yLr8oBCeK9RpaBnyIQ5yXAEFDERbH6xGjgyN76G3fNiG1azBH9ihdW0lKTyx68YD56FUYFL
h5ZpZr1eSWDy43vrq6qAd3q0BfJ+x0PaHpkVUgcn47CsYXfQUfJkE9okBvvHgKExwcfLedWspiBU
acOWM2KcRWgOTIexxW7EBPVmsGb1i0Dl5UYnDtYWdPeIVx2sClPJHI0udbmcMFbqrKhbizHFkZdb
TwchsPPzwnfE3TifUgq4EBs6z5iec8a1S51Z7CcXqtItYHQOkmu3KdJctKV9NFrzS360u3jUcaWT
dscqQX/JvlUbhaLAW5rjMvrJEn/qaZ66NAXLdd1nZiHYgYN/6HU9L2/XGL9Pc/ahcd2oSIh0/8mA
BjjtZC7HPQLJ1f9e2yXDLR81TzH3ciMpJE0AoXpn7lwOuYHUEEyzpM7dbgJ3e9fbPVyZNNO0mykZ
JZa7sL4CA1hr++vf0zFBE3EKgOdVuFD+JP8F66GWl9KWKS3ELGZIIYls3Z+jWD+i0O+I8smJFdqP
5H0VhFaYyTwtcMv90EOkf7++oWlZCLygnQJ3Er0EZvCO6iXIzQbo93wQP0QxxqhB+99TT07eVtFH
hK0A3o8ljl7mUeikoa/RQVzROaSSQUAuAVGqd7a13+V2YVuLLWsm44fyw604jVHep3njpoDybhWE
LAzGck6L/6rs34meN9HHgodXiznxxlfbm4cEzeDxLMdTj0d2fiPvYX/OlzbvSuYa77oFxgaLnY7k
+P5x78lsZ4hYqCFcqZkTj3T0IlJL7sB6viC6RoQLkin8iifMHdlS8qvflvPuhoYl4edpMduSHdgA
gweoxYoVQiekY0Kqkd+AQmEyGyeiVQVA+EU/pt0+H5P8sY0tJQk3Pdw73tTNbrJ6tonqeT5lIGTH
WqAQQ7JS5ptjLTikJ3f7z1NdAwxRYm+23lNFsDFygaSTCDxpMF5wsFaH2vxrUozddJ/RSs+g1usp
Woc6ulO8gevKEJxmZCV6QcP7W+RIUW3Hp6rlKYMtbHz1g9sFECWWYiQkghwM+NAlmFBLc/uGCk9/
Wu5BkqVOIvyptXXEBswZRTbUoeWrxatW5SHxEHt7YfUeMziSJSmh4pNOlQZP9xEm0VAOzqYa3aJL
m299emPyYE9zmDByRCHxAURfKv/wVTts2kct0lTB1hLvQVQebSwRIbY+opaq/44NYAv+zSK5L3PG
GzlX62YGbGyBSY4L0+svGlfOfHVgjHdc+385d4P1agIjzvz8kmKfMA2YrZjED62IOmqZBkWgiJfa
UMJQnC62ZgmESH/rb9DBGa/AYbL+7Yo97fkqAPTiRaHSf9PmtfrDEQIobUa3sYsbBwA2Zl+DvTpA
+QVNHJBamTQKZyQt+hPm3uc8wg4tz54tlF/IFq2VRI1PEjawVpcL/xKOBmTD7ZgnF5R6QDZWV8or
MRJTd2v1/vfR+ozgvLmJLMvBer04xLc5YBeBhow9wFyebC1NRs2G0S5eltk8BEC7HwJrJUY4bt9D
d4vlmfgHqKlSYRjyt3mUpqs7kecNpjMvw/xr2goWE4NMtGgwMUuSEXRqy+H5y1oj1euhTBOKRK6u
Mp7qcLKM9XIneHMj3gCTVmPO0xtDtwtu2mzuVATOAoIWEJI6Wh7szeeoaAPhiLJEhSU4qUyVoG7B
GPoCaj7JsNIbYR653P6schJoGT38Lplk+qVn0BkphDjHI7V81FzBY/FvWfKXe9Et72mnQqVKqWO2
CpIGbppES5cn2aU6akiPUAv0vNiK+cgK74uVAXK/xeli++oRsRdqTNUC0Ip8zXqQPiyD1kr50wzi
ARrhY2pgqLQkpmJp+aEPwFEXs0Ha58em/DaWdk5RDSTtHnc7pFkOZSKXL7I7fwz8eADJzeV01lhJ
c3egtoIf82dYGuS24a/anYxsAbnhX/k6uY0PZ6zlBDqWaBpsMB3s5ZECvXlfPn+4h8vGtPbsYisj
iamBaY1y/FFUw9Wjk78AiteZ7zTtTTUcb8NqqAy4d6CZu5Sh2Owb8YC3Fqae3qL3NR1foBaAzelK
x33Q3IaPgMp0Ib4aaaOUWI0WDR3+YO1bakSnzoWNRP/FIIq4odNcoIl5HwTPWDbNp6oJGNSW2PPL
GdRUFmP0i07Xh8N9/SOC1C7/JpHeOWLAlKaAAUPmndiVO8Olql5sBrYjRcC430uWx96KlXzE3jEp
rxpkSZnuLB9blFQAgl2q81uYvJW5RBmfyFMV1/hZHJWtllmOfiP4JljCQGK885I50LzuoK2wGc3d
2WhxLTm86M46pmIV9Hxw1/lAuaqzkORhdnJISGfd3SmnyaAAEpqvD+WHqxRYNuCdBfACLneQPQxt
XfPaITelLqoeRAXrOALW8bp5SEeq4uMVo0vlj8lkqI0f4COaI0sLxCKEWGHR3RJzGVSiaCzt/qtS
FksiAWfvZZ62kmaNWtuElSJ7qH+cd3W5rnYUA1yQ8PEXK7NuiseR8LRmlozip75PXMSJoww8TSyU
fk/DSoM1htFP6ajm4sTUC1fQ8stBcXtOpxgjQcklimwrgeSnwWkwSZWmOS0IG/4Nh77c7FU4y9Fs
P8zhxx0xhK2wpzMdPzPVFHEzRHRET6V8qSXok5Rs3v/bgSUmUG6I6gh4UIDcs5Nd8VpQ5vTDhLxK
o9/wbGh1KbBByw2ygf3eKFU5MGlTE6PsPxOh/41x4VJTyjRIszZWr9abfHzNh7JLo8eWK0SWpTLh
Q+1l+Ss8QXa3cab1ewaohOVlQxgpdIKklLIo0BkMbwstq2aAaFvQrwEFay9IWhntUQWbV6Bb5N8r
qfA886lJ9leJAWj05I+9xwAMhnH3zP1nrIrJN6sZGPtXQYYCzi8mKUTYgB1yqVtjylXacWaJHw8W
QNVc117J9/hQveKoWcma0R/70blJetnab47E4iAZxGpIwH0yHVFGvLphiIpyLeU5pweMh0r1f4ng
FghjvTa99BNcw2A0dvdLw+SVjpQ0StU/XoVXCpcGTon027a7KEOZJg0C97KY6H3XcTOyyro7HKiS
HhMk+htx6cd81DNhgCG8OjpiDnJIyWg2zHkQUS6yXeOpU2koeQUo0PUxLSidhfwsN6w8JP4FsfQn
fdlAdHEZO3lTLOOrlQykIbn4pt5HAwlUJVdpUS8SoyaymFlPMBUheHP2HTD45Zcw8CrhvoA/72ZK
dEyld6Wtg2PEz1uTI2cDPhkAYgBtTaSYiQVZPMxefUZIyWpGrNgfFVrNl6PuguqjT0yKXnpRLmJD
Yf9b1ZJEaewOD1tBLuF3eXSNPhW8E8U+7fiz9PUhi2NZD4rl9ThaOPydroKOvVA96LJfzG0XiR2I
qubQReBwUOxqvTO6b7zdZGmbBeY7zsDnyDKT6UqU9WazBLS/Cf63wM+4UoCw7x/yS1tRlDOjkNtL
jneE8dpCckxgTeybaWf+NGwqPtlTkeDs3y4kc5NTOKZWzf8tr2KPS4uexvLuPlGActjmfOD9HMxD
c+mUs+qWCgWAsXJiQqSZELgHU2QYz4ugX8lEXulZ15CRyD1IPyxbObtfddcQ7XEExhdOzPIXgu4R
XTxEybi5LqoSjuZaE/2RsgDH/tMW8uCOqm8OPa8cyjWNE6fDpRkAudvbgJGYWSO1wcco5j3dcqnm
XLqSqmg/fB/uQUt6BEI8C9jbpo2W64sFzaRAPhve09e+lLCM9B+05yto4+1WI+Ds35E+s5zMnund
w7nGr4lqw6XaHFhJ7xZUN1Ny5RWgaNOPlHxNvO3EvN0fWe0QxjwgeBTv23EpnTHSMlMfLBgEsQP7
J29qWvKitUH2JqfEbYImdlA8W85h5Qj9Yyb4ejkvurxLdqpuJe7DjpQcVjZOSHf4722GEGuI+nVU
1T2zKEBG1JMNJZAUFBHDqgVccB8XM1X+uAFPwqhAW9MkW2qskh7Yi4O7CxefHcOt3776SXyH2OFm
dpSvmVi4GssenYvTrVH8FpIDV+EU1/4F3uncADFX8aMGx3fYqD76saU73HdI+bxJm18beD57b3q3
PxlKONL2erPGNbbWNNY/zpNR1zqZuUavUSGtODd7WpElS6JCP6M9DFQwPfEIcI1Gf7+8HW7cetCv
AxFO39DJi79xomPlyR7XEZBSx8QX22PS7NQSKsC2L19UJB4QpraQRMryBSbJ4L1QGCTstiOouhwQ
q/5F5FofQFGI61EYwfWefG3BDoHRHJ+ZnX995om8LfX0MzZQBKoMKm+42WzhqTa5miqRhJwCmnbD
qA3QRgSZVlenA3krg29+RxFpMZN1RrJPKgpH8UpFfSawrYCgR2PdGQkNZHyBi+hRsxl8DvGvT5ow
vztvawyhrBB4dBaGjA1/IVfbEs4/14efAuwvdCgeb4ROxoLoBHEvrEFDDEPmm61gxUzfOmKEhj3D
VQYbsMKhqe3QOBnRg3tG5ZsijmsIW76oexT4HcRJfO+vQODzymtkZQ2UgLi18gH1UMbRpWR5rhh0
ZH9jIlyMCgIoZkJaMTiodv+6y6tK40IqU/YsoJ2Dadz9lFzz2pWA/bB2gd+Q3Dfz+LFHGCw8WOtQ
bxLY3dOrYjMTN6kWaiGMn8/2rHpcsaZ3JUycnwR/fJ3S4bdaklsMiYpQbDtHLfbnpjuApaGzYutm
RAVsJa0sl1DQMozO3Vokpu379J8IATtE7nFLTTk4PJ+1aTDOWsTUnZ/enQ2vVDzlf19cwggjokmE
+ajpCp9BmjAkLsmXwrWVs98SAuV0+MtQd+pNjXKdbGHhUYM32GVF1EHhvYeiB5EgwazIDRU5j0CG
OPyOf0ZnuhJU3yX1+1ds+Sw99zrpvivRj4rXwfXqvsagoMyaHmJQ55+NOWNud7q0iI+ByLM+1ozx
L813C03dMxQCCKT4GIyeRHprSW5rLIbR1nX30Ja9KToldq2yGc7kzmeyjhCFPlclEkiiN1I7e6/d
QuGofdFaEI5kMZ1IX5oSq7jPu4CuCCYP1e+qXRwkfiHUzuZbw0D6445ke11jGcILZGBJU1Ywyf6I
OLKU0g6gynSoN/TsJmyjVeVSN7Io2la9hnjdM/Va4Ll4SJ3p15YwiiCIEWoX31PMeAsrUA4atWll
Kuyvyprq/0O1pjlNgJIcdO/obL1x2xRU7j4kRs4gx6UlfvoFZOT3jbseYFkDtid7YV5OjcRAghA+
j+x9KOUIstPTqoFoDgCrmBoz236PaUjGd6exYlOzsxJ6a8qNJX8he7qwn1MuXbcITDQCxRvz9vel
jJ0wWoLoutPYsRUcXbHiELJFIyUSitxn5ZFmyneKKJpeeInBgv3rKBHVmp/Z1/YY8YTUeeDJUGI+
6UVexeOkvjvyoaJ/3D8j188d8xfy31j0eBNoVFr2ZU6rm9s6QtB3Hb4mnEvVHkXLLp5vMrNaN3nq
YdO88PPwnJqUBHnIcJYBWnvJjegijfgRri4vDHKpFApyC6w4njX1DWHvrpeAr+HJC3qiRbszcuEN
BRHwRoiAXWGKAYsAQOgCKncOw6xYDQuHLqk9967HnF45bJwbFG4yvXPi7QFlRe8JWHS9pmJalrQk
7hxyADJQaeZekGSrsz34SJS0BVfXXrfsgrvh2nWGK0hkTee9szfje073Mral0B/OlmluS7l7GgAK
NdXwoFlRsQVPd6gqj7s2oiUNsvDFfJEl5Ts12Qr+CsXRqUr0a9bnWiSyEy1TyTwFRsMKaElg+sGs
nytEgE9n5zuTNYMaW0BGDn8q1zc01xJEyku2Lob4EWPmaVhnXWJV3+g5NGziJuPRTVMz/80CMKd2
vothytBc5QqlakwNPiU7ROFfTjsAO9LllzeRpLQXotwI4Rt8PoWOzq9fY4HFO5GZHyW6F5L04Uyx
BE5bNl4XXLr9PzNhnY+EW98zWy75qb5RG2pwjt53f/NI+2Y9aeTNPjfAo29DU5qZ78Gv2Bqn7x2p
ZSoDyrgKICqkwwfuaqpl1W94KyXxhbEur/aQD5bsR/Zt/GTBHdFwU8tisCAMIyzPtzrSrw+E5Qmn
98CrQ62hfRO/99TE/+SFL4Oze70HGL8bJ1suydvAu3dKWAF02IimO8bl49kzEU09Zw/DifK/uBu6
iNr2Ca/+JBEhbdt3DO1xQkwJoOfZbBea01oLNx/58UWfcWgs9mxcULzjC9Dk6LQ/eeHnB98rgWR0
+GZNnEI3kZSi0Gp6gFVhASx5USvT9kzqtkJ/9dHG2pbyTMSPfhGg3Z6smqoVShPll12VCAPTRo1Q
5ICKU2SxBX9MH8zXJ/nIfCH4Z2xTr3w+Cs6lLVmbb3YuVlG4EWjsMEdCW0qVH2o4T3RzMNUZiXN0
DkhBbhERXaxeZ5GwZbWN4ILd3dC6f4FyopmIU1kPeLjKJ5WX0juEDZCWUg6440LJHPxKeAWlewO5
ppuaQViNHvMzgPBOp1fF5TAjviC4Un0uJ5k2PhFFLv1mMBH6yQytzPzfNyxJ1neBBqPIJCapqCOY
BCx4K4iuFNhGB6tMF89P4h7Z6IK4z6LQtVX0EfYtQ9MIBdTpqYaSjFyP5tG5S4Hh0OcYE5SEW4B8
zMRziw0XNofgcfDui03FiOrsxbkjqSN605bYUnezZ0PEB4Vh8sJyRClVFw53Q6FPxZVPMdnMNSH9
yiwXK8pxpUxMC+GUFqfpUFNavAMU27TGYvhD1Ta7LaPpv2HL17T2XbEsJBIUC8+o4EhqYfCBWFo6
jBMAIub2MPOEf+f2WTtrtf/MBpLzrYb/C/RlEyXoqhB0MTqqwwx116blDiF/gEMVAwHuZc5E2ZHj
i9UBZMFfyektA2uNM1Zwj8wcKrRWdvhFq707zEztQkSjdN+r7btaxt32oYApfBlw7hkb9e0fYf7+
OlOSOHngsqB5rju7749k9yfgs0RiULsZyR5O5mtucsHSxVlDz/gp4+QU3u3AgmjOXBEsp+dNKX63
wU5qusgNV4s1McactiVP0QrEXBchyhi9LLoRtNlaImOaDH82L296OQYLZUyV2NT7LfLy2/hwiJAd
idgpnjejhB46MDr00gQ6p43+5ZBkFOzorXBULoQwgVMNV253T3BqtsqPeG4bpk9B734/K6Ycz9LQ
M4tEznwxqcVehcPjmBZoKM2/KsYeuIMCi0vQXhets+1HFmsTIAzhTfPTV6LI8EYRkFJtLjujJvGr
eRkNtHlx30YNCYvl7UYHr1Upu18Z5zAozvMUGem7nDeISVdN1NwepKV2Op3ohTdw/WleqQeYLzUG
LNd4ZiZA+n5Gob2vP7ixEhqX7C7QeD0xe5+ueh+IWCSphDWA1gOn5ag7ku/KB0eSAbx+tIMwj4dy
zm4Pp23elAfhAb6yLlcxYzLVhYn/1cxVD6DQxn7joLUQgGAn9jgWJ+fpiDVFzNzSeCIwR/f9ZI+y
rkbAg3Y8BHUhyOG39sbIga+R2eeWOa2GmYsI08BI82IbuOJ7W96mclPFUZEQEeDGIZgh4jUHOvlk
ePArNW0diUNhz0gnQgXvi4fyad2kBWziWB+5ckwJ4wosvyHiVwB+uyjPK6m/dznRF6rK3kdzt/mv
tlIzr5z4Bwa7/LADm/mTSlBIaAVxUxD7k/dxIngf/krL8F/Jxqm1yTqBEBAx+UCCXmAxILyjUW4U
e7d2YRobQ5KMJCFGxhmlvl0uv59ds3E8C5QQcvDNw64uYtGZ/aC/lPwFfZXfqIwLnAtCy17nU+Dc
TBYmxtsbTKTxMjnMvNBD/wTT6lSWIqU0aSL+5edctboIi9LRR4MU9Fi4ytuA9oVrGxpg8ZkZDG+V
EQGTprBR5Itg1d0NJbTnYMjdFkeEAqdxxJ/7jP7Ics5XE2rdkMSO8JOrK7IzZKJVLQYSAHDPmasK
b+9okZTAqMoD5CCa8D2ik2EL1r6ihK3dGBbsvjLJYHKYVZYmxd7H5X1VLm/fp3ufXAFzKzLkNxzl
VXs0rYDY2XyuvUhNUeNObvK8LcwnpgHWQiOisHT3hKXRSyaSIbfpOyjDV5r1B53DAg/rIND8gGSY
FJpwdraNv9+WQhw7QrHE3UAEAQofE1BFtIP5ua+KP+EcZYD74uVVyldggFSSoA8J0amP69JNIqyc
Ww1c8PsojtFZm7bzLgzBlURO1sgKg/Nw8jQAT7oGSEFTzEIwTlswW19oIggGvxA5PJzvfrPfTHd8
CxYMFpWNJ0K9GEm5zJrlNK+zBcw17UYye+J1+Gj0c7WHwxFdQOBY2Ou/RQZtqpXDjYMcXgTIvD1m
HBfL5vZvIf+jsGF1k1QCDBpr5WX9nz/9XCsjsOfxJgbQR+y+2inXiJTKiHNiUcolxMlAj4U8gWYW
RTQrRn2LLG9vAn+KoxniSPTyls840WjB/HJyyNB0/2/7UPeh+7NSKatJ6Eg4o0hce7j9VBSbraaG
N5oBmJOxJfd6WQRDS/wcZFL3hhT/ElTzxBuQI/prhIwu3H+uv5LmMTm6zV+m3kWNdrWyCrYO6Hjr
146RLZbL9oQF1sL43iwIfxqszcgfoBOO5JjKxoGijEoIVRftRQ4xnYi4PEG/Xsewx5mQvr9PiNp5
3HGy50eIjlZt++N75b1XxVVuRJ2yLMlS/s40hlRX51sWr8Gs1nGzBg24dXPeZuOG2rgXpcY7Fokp
Gjml2MmeYydZHj9U64xmCJ+hfU9roJ6KgMkYaVamDdhwiptfRiytBtx3btqOjOhD2hP243fepVb+
AOgJC4qxZgjxCBktwdYTx3l/as3gulHXgM8KSa0bIuuU65OLYuSVCWL5mhnclR/UB9URfq/PhL5s
XzHRIIz3ns4rIh9LkoYhdwKZfNMRgOYixKT5/8LhZJjbgsvh6jDwiy1InoU90ks6P4lqcGA1UVH5
vTzfBVsm5JxluYvJBxiv59ae/awNfOWFLQFKCbaWeUa+OSSp2RIPKBMM+clWLm6vZxSHTBoERZYp
YXaM44yBsiMc21KhvKPx7TXxqH2rZUnt/gG84vtjvdyCDCT0D5FvOYBbfCH/aJG4b4cXW1/g6fQl
z12z16z8QTg4yEJuhTv7T9nLVeDLG1BbFIwGSr8X+3fVm1YOBquD2VHK4MscL3Tj9y+ALqsjsszM
0Zjr9m+mRZNhu+TYWZKVCEy1YJBSJ2EOiGkKhBJz+U0KGUuuNqNPzZfjOsnLhdveWmnZLbI2c1eZ
6RkWTVt1td86ER53RYjNinRjrLBlBhfzuL5inLfR0JxQuuSXxRg+XBigY60r1J+QQ1TzluQIrABg
T3rwIGQy2jHo0RzFPpm2QNwDSxODvzqbxcbc3kNEwt5bbsdSkJ5jLx+xARxE260oCyNAOOyRTEpH
PbqHTIYEXvKjLZFA6K/MCTzGRvqE1xicsfPMVVEtg8sojxqe7GICAFGDB1+tgteicCSbqguxH8cm
FlO4AqoAhbrsagpFhnakR5AbgFVYLxr3Mm9NyJwm/4PgAmtjmTUA7uB1Z2DfxVKw0bK6f4mNN1zc
o256Mp1MnAVU4yLXj9/IhSeLAh8eDuJh5omkJZTVNIvm9YEEtbd3K+yNA3eINOcBHIyQgttEwnUm
wpH/x7q7k4Wmf+8V6tQLukGOVAq4E8YgBN9gFR3xeGBfY30WzBcta3NcuYYYEfZDQ9GO+JWZTthS
xKKJsVyURlHbcehcLIWS/nZwEYTdzrjTaGzn24LfomKRzbhpv7uZEIKUn1drCqR+j8gaXwI32tFt
ozFAigjU+OUCWrFBwUM5FadZx8wJ0UqtnPiylLrdpi7dBZADtNqCH3vYafBHX+WKDNf+n9/s7qFR
RRGb+UeP0tlqB6bpFPBmJBdda19f5h0cqkZBlAfpBAJY6KAIO2idMzFjZXYwmQvqdsKtvlZJ2xT3
H+VJ0NM04sLPE4y4Asf9sNzbHEyg+ASj8JLRODM6JCD3WhekQ7lHMU5OHQMx8wlM/Z9796M3xmf4
xxa+k3mE5dTXdC1FxcpTnbQGW9I+0qHgBXMzlc16Rs1s6muj4PXNA4nHptiOddfFdZ+xyVQikKFE
0CGKqopX3WTksccOVV4tDVgAg068XNnhVghfW21zbL/SvyJs2Q/Gmznx0cXvwGCLBuuB4PKFJ2p8
/MjO+LCYZK5/PY5WEKOgpdtOE/L3nj71NSPHz6OQT/E5xszYioKf21CHRB+Gl4TAEMLnU113Ipu7
Y0zggqtMxWejfCIZpxzJehMtqQeNZAaMuAoG+kyKxvjjUaD4NTMsHdamc/wA7UpwTGijwuC5tVyt
eyOnEAKBVn7bnkptX2pg0hI3rIC7TuAeNFr81xIu23mpabkmDDn1BqKFWjUqnLWv4ecRxeNkGcHI
0XITaOPNSa7wEPKh1w2TqG25jX+fizGtSK/Jvm161mK1k0Ndugmu4YogqF5qM1QIgQTYu5d0RgIV
BWT9oXEnWHrHiH5Jnl+4UIVbSQl0eu/lijvwpCYztxquKmQHNk3/rmhPQvrHwYKh7aPh3X05/zqc
ZSJsHyA6QOOutiSBw72kT8VrHI8Vi14AlU5hyOhSeRm9LdRzFSH/64l51vxMjZkN/fw+Q/LhD8sQ
ksr/M0CoYhxNzrZyZSLAnH7pX/JlCpCV8GNWpDfmFsL32FlJfj9buy2dln8dGJuqbKD5Vqb1NAeg
ww7tv9Ek7sL48t/P2ibUmt94EpN95tAlneFqCAdZxDNghdFNUffbhakApucgLtBF7lg6QLT/t8Xe
GqgtE1BgebwwRrifKNVxKhXT37vtubJujLgW7FUFRZ80xCSdtacg3lFDxmnYLyMi2WxfgdE6wxzE
jpvENQ8Yc/12aT5/BGOcdNsLwc4echuvmp/8bBEuf8FT/mRd+w1PZNMIlEaiOlemXGHsX0SyFq5/
yAyFjA/OQaT31LMVX1vosRPYGlALlfGvNKfsY3ngAVueMgA/mhX98vtwtpSJL/6V0knJ0nW33BAU
GAhTl6MHbrJIW7ZJorMd6eSW7q43OQmopjpK6ceop39XCGFnDXfBknS2z9LcJSohBH725cAPWxLq
6h2eRIcczJLbVQzDzcwwZzFKHAORaeUadqRFPtK6NmsMt50WFTjhdruig07/1gfH82WxNazaTp0P
bG20smZPH8JH3wOkavPGSoWD0NewKpXaVDV8v1fkOP/+lFVWFqxaiZ1hrf7YlLJAlmqvD4EJFmk1
V12QynYL4+Nm8M+0uzaeE4IPWW3oc9ZbdeqeoqXEEd0qdhB2lh50O/sRjMiF1Y+dHHiym77zoqkK
c4+U7V4XV/CibgHCcQ7NKzW4ZyGvzkbyKx5pSGzE1+6h1gNSv1s7a/QHimaG/C+g7/h3q6o8dMUV
9Ytg6uohJx7TeHfsoR89ZKL6vOQevy8tzsO0a8/dExTxMM4DM8KI9XzRi2ClC7Op9RD/ZQaBUraX
tQ6wHutdvumEbXJJcaOaRh3K4diJGS7iUNlFRkCQbt4T+iGljxEZr/tigVutkzrXI3GGS0H4lLqo
shAz6hNqDEuenpMku+jSLd4SF4OADFQedOae1ad0PGJUQvBhnTMI83v4In3ryo28McHy7PHeL3xh
XKne3lgfe+wSzCrrp9qRZHfRKZYsuy9hvsrTBx/6z9kv0niuGb5x3IOwZn8Rk5l3GuKyUGe4EvX1
S8DgnOtT1YxDSsNN1/EDq5nH0rfQan5Iu02LO1rqfcGwypyruoO+CsPJoFauM4Y0eskhMNJum/qv
DbgvoQ5w+sRdK8jcLAlstfQXxKYh5oToiH2pZwDM1S7o09vsUzFIYU9F+uPf2GYFLOJjdz+e6IJ4
+QiRERRribFPVq+bbKSvZGSilXsCbxPKtYwvm/sazjL9EHXag17EaZq93S58JneRZW9AOOGbfutD
5qZkrdZtydwYJS3ivxXn36UFwhuxPsRIMTOCfep0QaM8VAsnH2bZmk/JU7Pn2UDQ/cwvkM4twWUo
AOad1JFnvP5l+sqXyB+IQaz6rfe6PPt9E4mZwX60DdGixtL5dQXPdjtEUA/EgRN5dNQsrlJM8DWF
oS7jZWU55Junj/+ZGyK4q8k1EnogoYGDTGpVR0KgGHXnOHFf68XH4Zw1QNHOKyg1L9I+34GcCMin
eShYOCHazozLpSOUBJbIGvwj1XiI7tXQZYIAPUxaa/2s47MnXJaHDCMeS3Fdq26TOGQtglfYymKt
gXSEVMM1UGwNZlOL/PGMOYD88yflA/BM0xlv7UH2BQfoIXxykqb5ZJGGy+J12ynYyBt3e1SjP99Z
V6nwlFU8/e/9h3krxnpwbx8mT0GaGMu5GtwbiwYgjSg22YNL6n8KarpCiucb0QFktrHJQEg6BdkA
FvaC8waLf2+AaRV7ltGxb3ih9YrVvPh7159YrjvE2cq03uB/HuyGQMhVkaFsErUmdoiole4yXikA
x74/l+DK5YUtJvay0hdKT9EF5GWrkDY6FaorlpiUqBOO9wAV300NaEvRsulZQ103kKyZVz+lWfpz
B7gtSdqy7GQKpcq8lchUe7W2L07QBDC1HFFAqX+RQutRHt2jrc6toeIHHDTi/N3cQXCoEAv8TZUr
7zfy8QQwylC0D21P02QJmaGz8ClA1GyHDG+IsvdTLNHVNM5U2L4kiWNK7wfaHE9IoTvdqI3+sTTa
A1QA1R432lNtuiKJ446DO5XxpwgjtdfWxwaHdLWYAsBaYJOUM+w/we/p1CKlX8QD1xqqJWu7LgQI
UJjhfdl8wLMYZO0t/LiNmJ0uDTzSscD/KtB45kvJBHQW1LwihELuTZu699NJ0FYo2SvSwzshJnWK
USnXsHtJ40nvaYMW673pV6JizU4/s2QLYDVaARehKVydSSXGWWYraprzRR3J6ICY8htRQiBIAws/
674L2xqwHDeeFpQ+uJCNElh6Qe6KcK7JJ7gi5oa0xPK6iFJEKEjIZzvdDLGp514wVX1++YuSHeBU
kWjpS9aRXUguB6dUcdOKfYm1JxKIgmsxUzBsOLV4VGxsVuX7VGObZ4To2IKm0SQsVYK3ZjsXu9fs
XmQxOoizpvXIJBJ+xuFqVI4Jtl3j1j58jBDx5Q2oCnbxHgEmUJPo5PFrMYhR5SG0BI+MV355qhG3
rwhfoFRMyyuTvHlmTMZaV1KaKwLHaBQ9txaOEWnxW0iBWcv0LPlbZU+DSNuJKlr4SXSjh80dKRfp
5ASTW20yFwYKErRF2Yj6kNaVjdERa+XET2gPBYXReWowmj2VnSwVpgnzGUXyOSWv6Aaf8oexNEUJ
hYm4Qe9gmxQyJdFnO7eey28P/7DcFbiKfZer++cURtz5QMfayvDZclOMErtQdC1o+R44d13Anf2j
Oazydyw2+xkTtbsAQMdcgrtB96jOwGB+Mg1Fdgty/XQdWgNvBy0+i/GFNwGlKSZfljhiN97HGh27
2j9ZAmlUpGZE90dkdrbA7BCXoy9H9LrMOia9+M45SFgzwvTZhZvKXdsZJVYptVtC73zLW6zJfydd
UhciscjaUL6TH14+koRmMXTRWSy7zPcy2gUMdY1lavsD5JUzzSPC7X30KDnfSkClrRF0Bazg4vEW
/RP1PJFrKkjRDKV6vKwLE1NXkaSYhb+zEuX+CJFev5DHv+1nsSPoBM+TPppRV6cPmDpDixss0q8l
FBIM1aUlbwhYshfzdNDqMI7Vm4HGG3fvHrcjnk69RO7MCRO2HmzFPdxdwdgEKsEHuT+UR5fCpKyY
6Xttb01U7EmOChwur9wsw52lVYAFSFg1sdOWZty4/UoYnJ+1QGBwTeu/jDVUc3KVcwqszOPCcVl8
ALNkBL4Czx0W+Sr0A3TkY2G+gegBRyHERNRYO2q6gF+L4cikRjC5fc1UWTO7aon9DOFG0ihPqK8O
z37eicOIeICXAK/1yEsum7Mu8G5NUXopVRIArPv3Zc4moEpiehlljYFb7J20xGC6yrSSvrDNA59y
F3kahy0rwxvr8O15hHTfnX1Yn57GAJeqs6hdZf1IdiT+g+QM/ojNAa/d/3EG+wakht2a5c43vyOs
q9NG+sr9FeUp7W7wZYeRAs0x8iBvFYSBx79IFLofzgeeU1tF/EcIdVU6POWIC6/JF0eKKysb5TLX
njv3hU8CPEoIdx+WSyizRnKePYcRIBEJT1hgVdKYw79HPsPAtnBdF+jM9nP1Gl9gs5WbKDLT36qc
FscUwcsrngVsSCtnOlwW1yYFD8CL+quMHzdlFe0XuLRl/n8gW7Oem6XBjVwgYgpRFUdztUemBBXD
g1EJWgmZYD/Ub4nWflBtA3I768re6QY6XHOx/Gs7XchcB6N1PlBeySr09p7sKvSo87GQsOEpipzK
BXBBQw1H5IW99v+totMR1LIftAvVKSQokcP5C51FnTPK/UCvcB4fO34U74Zd6NZXcS8nELM/Rtlv
OTlmtpzrn4c/v0XDZ0hXBoX+vzEL96KQE41Ev7VseYVGxLqZNtWGinJAc7FM/sv328VOac95kjg1
tHLfMImIH+WTVgojfyLHjcTFs4A7NkbUsZgXK9Z3n83E2cq0sYkpZgC4I0L13e59ihsoZNNde8aa
Q4Z5QbDuOJ0Ti2gl1Q9+6RzMc4xfEw0bpu2FNlipzt9NhbsapMPtxN3sjFgh3JlS9+Fo2rCi/4Tm
BAVb+m/t94Ez2erh9pPdCA+SvgXIaJZOvTWPvjhiWBHj5YHBb85PfleYzNvWmbzHD2J7+Y5zztjp
HMa8s0xZ9+4TQvCC/CKN8nt2TiJMZK+eoeXeSDYpzPQI4Puv1nLmPYE3MPKeMA9dSaJpNfOJAB6d
PeJTsDxG6FQy8g1sop0YLDMrgKwG+afj8rAMlBqUf4UT+e72QqSk+C13Tq8mmg/jpv+GYkBL0T01
s3rstiOuSsGofYVhxQwncUDmOFVzUbkv3BeRU/+R5UmoHQmGx/z1QE0hCa6Bokgi3WCFo1iVhujy
NasAfvHInNlH6Qov+g1n2SzEn0DRn0+R5X6tFasl5kyrCfsJKtPl3UOQHGs1YaH0BPRQCqRNGaqm
NKBjKgKxv8usnueVA9oh80X+f21RTn0hqQHSZX2BPKZBTnpin+dXh64edqal6JB6jc8SAW4DO8uK
hQNe1wTUrxEVkfNo0LyZC4iY8oc1gvg9iCHjPEH0ES7nlj5Esi3z/cLm0rXZ8XTdbShNHC2qzpaS
LcXQapOGFvJkdlk2V495v25XTgKsXXxW0NQVxOclOA1RTDNxgbdGUjqO2iikHhdHGCBsq7eJSbtX
0HkFad6kJSsx6NJY4+5uvT4Ei9/IgGnQOvKvs0xzykkfMxjczynypvljltLwEPcnhineIjs0vZCO
KssIQ9unTU677zhXTRt6TM2Py1j4LGwi5/gO1RamDEi1Y1lk6X0dQf1VeEb8hkjTdPDGUxjQPXLx
naHqxtu3RRV1tytU9jqEPh9zThqaANNrLjolV/YgiisnfA/6TD691VsmTINN39bnmAUMpbKVZINO
G0DSfj/IiFdml2QwSso/CKFfvk4GgOi1N7CMmtERe0sDDnn9MGgI8qTuWX1MjL1LqwsoP9qMInvQ
D4vC8rMj8gvKQ+ZfZeJ44dlE7bAHTtnyA/k9zwgV2loA65Dn5DUq/5ZJkMndg3o8Yc/xhw2exRwS
9FhwJG9zEmLn5tX/OLjFCb6Afo6erTvQiOYnIPYjjNbJL+5IDVKCVmV+9Rgu4Pj27UETDNOGoJMx
UrYzD0lie6RkuPQJ3bnQ0b9PhCoPsCiN6sx0pZ52uhXxqlTkvHHx3WSiW9EQCO1KOnv8cbbdPJpA
l9xuM6/nerB9/NQfXotMg/svFaAwKR3wHxTma+v+7rBwIGLxCFdS1NgdAgfvNnL/a4+3D/PHo1HQ
TTjT9Q70rzmqVoOxuHb4eswRfpJ4dAcKgnZKUB1t6l+yDSx9y9GMulh9CK+kZecuSh1tELafBtO7
IKBRhRpURfQJIrhD2p+/EbJe5r3P964/dCqMpaZI1w6ssI/iIhbRZB7TTxeDat7XXP1Pj2/E/NIb
IAeZDIWWrqfN36YDbiXVHbiZnLWw6r/YBhZ8G1VbXwLC1DGd2CVqGmmansk8HhUj8qMgGP3RDR7L
sILsZ0PXE7vuGW81aGzO5JllEY3ggErPyOfrgxflfbJobdT3EcT6O8+0iAwciYlavFE681KKpEg+
dOySSbjI+HY4/60xZs6Dl8Tna81SEq95uOSJmmpw5fi83tvaAi7o98ThnPwCpguYCwWf39onv6rf
a8HGiZ0OiTy1fSvn7bKjj2Adg4gJ+Aoi6y7Bw6XKm57jaeIHVFo1BB3KPtpcRkDPoVaBDeJVI+BR
o9c+qnSiXtLQJuA6aH5TBDPh9vNE0vTzHxwdhiGsIl2hv9zKxTgh1tRhMIYg4Vr0AKFguQOjzv6l
QDkJXZlpdnYdu8sFRio3Wm7u/CJU7aOR7+nrzZ4sRKo2EJ53IRZMe1nt2MCDw6mS1FhjywsOcDmP
24IVW9DjciU4C/+DN4d8AW53TleurhUmO3Md/Kc0lOQi8Csn74bnnDv5vywoqNPTM4NjfqYiafac
Z+vorSiz4XlC2MO+bOm3m/feRr9yD/iRwotAgbANp2hJThlz1hYgtH94Bhz+O3Tt+CcSzu6kx8VS
at9B7r/7ZM506QFKgfLQEMuaeofWxU7C+yR6BCPThuw1Q4fttB4dLfLzDH/FlDVpYjwu43wV22jo
l55zs/AuRIR7UNDCdjn60INZk71SmpJedYbQh1f3NWC4R5CKSh2mgKYdeU72+w6GuqJkTWRecPMa
pdQ/fdWBBLJnFYQUVvASM3fvF5HnmizhDVhWPofd+P9cHg77sRWURzl/+mzVA+kdTXRvPKEBPgR7
7WmKVzZn99MHRMrzmviX0ogP1QBDjso6nQ1ffP9qGZSKt2b4xx9lGpOweIGIQ/USP2QIodSlbxo8
e/ZfcfohuKWytkuTdKxpZ5QPMAy+gBp7tNgM0c9UMgtT0oLSigf/z+HnRQ8l/rSPQ9cwi+NfADOr
NDT8zqgyISMtO9MldmIKSR80SJaS76UakBfqEitaQ2PdpBd5dIaIlxwpBAzhv/xDj0KWpcCqpJkv
cR+ttogUGwE4S7braXdEZY/jx2LC5uaM/5XN0vEq89nJ+8tEUELTxxfDiv2Sat/A4WtW4+/La0hX
s23zSv7MuCLyk5uV7K7vPBnCABNFhUqj8ATpJd1h1k1XLbJd/gQ+G9UWt4eg4pPt+Zpfd3P+0G9M
jGIN2gfRPRUIR3v2wxdIw6vWxPV/HvePbf5/gu4aR6yHvHWdtrG2wa7x43ZKWrRGMuA+yTIpHamX
IWVLl9HZOieOW8gmO2325zgyHqVp7N2wZorneOrfsEfbyBKSXEg0EdXFrYw1QiRjz4Mc3oRVh59Q
Wx7X6Te1Fvur1VFWdJG+TJc9hxv/cODxYOuok8NCtv67jM4bkwjAgfKjMlB0veXwAZ4udNTaUMCo
JUsOKrkC9DsC5U/fUd8O0iNmA9u4856ej2lSgIPPAGUWLOudLLG4z/ss+OpvC5BQ/aWLRU8CmmIO
7OVzxChCRgxQFly/eadeqUVcVJ30lmIJsumot49xzTalaQS03+2p+afHdpuJDZcsppvw+It6th/c
gtPU8utmqiLHszLW34ySCgTBGhENL0NsfwP30R/Ns7N6DJCLst8xZhN2lWaLjXQPRmpUjfMpYmRb
Shx38oDIkrpasmvdVqBeK166kJ2SpDyF+HkRK5LtP4HWyVrSztNwI0mvQkQRpKvZd401iAMOMq7H
k6OxhX/wyOt47AIiMgozZ1J8kDccGJgsu1i4A3LXvMmYfwKPssyIaohl4hbKN4dHPLS57wPu9gmw
naSI7DNyKWDfcMQ+n4/6ZvYkcDKp9nWL/BdtCWA0eojHKdY0elhTIBekchdbD0KoN7yYV8zbpfXr
VjbhWqeybxMnleTuf4WbOAp3r5QwTSiiDsd/cYQsJh9xg+xuxsH6agM0GHBGywyB+mh+SLydL9nr
9auR4bu7py2o/I+IShorzIDpmosDjQtCbwVSNCbLE8jDd38dw9OGJAWRMhlZKtp/VeoKSFArrA5z
QnBngVJZ9vxOjoCgEuVGGwfdA6/1dD/g5FwNGY9mNkCPTMif4Ui7knlMfp1maXZswOrePUuFM1tk
pIMPOmYR3QcdR6/UeVtfK6y9x/q4VHII68X9a+nVZQIcGEXgkyEA50NlUcWI/PYAhs5Np0GF6JeK
7Iz9Z3PxkFs9bgEemyGDrWyNcCJrXrpp1Q0iBY3PQgU9j/soTir06NeJvvHf8ByhDEzM8rwgkTKo
tQSYNqTTZGd7oFWNIttsfGlvZ3AkjTKGyf9xftzVKqFIgSQcT1rh0B0HSx1eNDyGsR3fuqCHZl/e
YU+NOrPK44v+22QzvtPyilpQ07eytNJRfTsEbwDvqmYMLPV4YkvukP2QrglCirzle8nme5HQCNFW
c5zbffqQUbrrM506jFALDbcmSYaikCVhLi7TjvKpSFIPYHYByXgmRf2kMbfdnLuIl11WKShYh2VN
e2DV6EpJEu9E8UFuk4pUQCYrDf835vkMJEn6dbjB3ZZS8IBc+mR7SHcsDpYCOg1ehSnm6j246LmT
QrfX3Gk0LRYfBFgjKr5yrRCAUZFP8bM9FgVmSo0ha/MNVB1zmjYazpJa14fKM0ulOplJt6c1YSAN
pL6krfJhER8fuaN6PpZAe7uNOCMk1Vay5doFB84o5blNbtMCesw0d+ETJHuu4YhdBj4Xk5eVst09
wEyEqrwL1UuduCKi0ePBJMDeCX0NwePwKP3jARKaQkExBmdCcMdmGDy6pf89yG7NsWkMPfLSwTHW
MF8t58HWGbkezfQRhHKVTF7ZXhLtkij/3iXM8xpjv1bk9moLLgJgp/6Dm83fUCCnk/U3RDTZI7Jb
GKSoO4My6hV8m/bMbMIfu/1aVI3Etf1SY7yt4NGexbYZz2bmYrjLPYu4U9YWvnLrNWjLoirFNnR1
a8zYVqoVa8QvO+U8U+bFXEFiD5T8+5WuJFRt2N0EVeXqk6QHL6NvnR5yOpBJZKwifPXebSh4pvEN
jgbxLj0HHLLsFn+sl+hZoX0W+LUlzO6eqng2yZTeEfIWiXegmyVpnFQqjcuIhdqRNpPAPple/Kbe
XqsWh597PtgFPm48uLqd67/dNgJBedJTVuteenJjbMS6r2VbPCA68MRwBB0MTIsVOGIbVFQgvfC9
P/aJ5IJaSbjUetJUEHH7RRXwUL+XCCB2sV36Us3Bzi5FWxx8ma9Vz2dMBSXNpZ5MdZoxcrFZlMV1
XXc+jD7kudt3As0EGK0rCCCFbMQ19YzVxfGeAoc910gO60b3C7LDYmg53CCZitx5N/+fMgko2Aij
N//92NPHEpaSB7adFqU5VztfkhawauQWnsFByDdD1emASTG/dkQKOMvIrLfTQIriuD3o3mWUBVB/
bch8Q4BD1hnOTflkYxBhtticQRlaUZz+UyI1Skng+i6DfRkCFkPQdcw7bjayVQ4me/H7y6Z+UKJj
VFDYM7s8wLleVl/KL59wOimr1Du/e/WcUAXbNX66UVLA/lItodwArAou51SVLxoCt0jQUckdoytT
PdTywHpVFbia9q5WCa6fCdPrsA4o8Pf9Tmr6An2PSUEgA1KoUek72zZMYD3GTDiiSuOy4hkU9m2d
Ucba71oYk8RGKOM+XAeoce+Dqi7JCMZ+cwQ0d4mLzv3DdD6ZVfTHN5cKA+1vGdvMjHREG5sd9Gbs
LSURThTo8t8r0ybovCi/8iO9X6ncHPso8sYoDN8UnzepDTTU3bixCN8anR1nRRwmn5cpFVop5c6g
et70AVUg2tdKwmRtk+YidhkJVmNAgB8CgVvRqoe75qJ5b4GMFYnnc1cCUwfYxZObmh/OSNufXvyF
JfO/sOvR6vtT8G1xpSeIVhMIwvcTrT/nr71XnmSmep2RnMfJ8CpP9gf5nH0xI1A5rRohiSxre2hx
t0BH632hpXKdEmzMfjbXZHoDSnsTw44yYr+wznWtVaDrmnXPga7cvegxFEJzWj4yJGApE6WSX+2p
HtWatH27pAEezVGnQMsyhVe0FgR26EGrtXDDN1iQqsalso0WZGh7TOkUJpfTvgOAyGYC2fYLboI9
iqkroDR4LxZU+iknMRGo0WdjNYtWthDsfNJPW2YgbOTvUMhWC7NXevxWU4wyxHYaUvkOWCPuWLJ/
E4Zwvjy/w2Wc8OdxhEiZkqMHiTejoO0Gj0nYTd/nRTSj6L14NeYMLPWAUWjWVxaU716l0XfE47zZ
Mc7CJA8/deIXDWEeKpvL5+EWOCyFMeSraQQirtW1BqAAOw+XWqA7FR6BpvJ9yQT4Xgto2mFbUEHE
iPODVqbgQ1U7Pfucop/e5V8ST4lSmDXvd0gumqtnqwTrD7l2rGr0soKxSzQKdLbWlC50ltp6b7yF
W8aFoeXkELAU2BE7mBZHagD3f38RYn69mqyKfb1fKqv2wLA1tLgyXsT55qPoYmiOIv/fs6lg8M8+
o/EIbB8FBuZQn30/TG/ZPb9DYVCH0cP3xPfNdfQ4Pha6RO/7DrxaPEefwATfSSx5+1cBm5qI1kfC
tjGDx3d9eUvOTeu/7H3IMZOosoKUdq/8Rw8BzDTlqwNcXBgqWLpWfOcHy+PWFke32uY+j6dP8zOX
XL6hmlRKQ6Faj01wjmTq8RdaaSxrn1X/wFpVqPpYWozmdcOL+cirZtZ50U8hgfLoR0HuEVosi2Zc
aAbMJUZYDt7GhQFkBMpfSD/gtDAgL9e8YK1x9X+hH0QfYDkV1cGJGlaVPd+kchttRYzT31hCMKMm
cHXqgPnizyURIRMzT4cC7j3xf2xUWEr4ETf1LgRPKcTZwgo1WEdVfESSygfLdc0BuZxdh20UpHcx
sOGvn5A6xbltu6YaHTKX+A6Dd0AcW22ryu8O431dPFdzKvUqfg41272walygL7PGbeB5jhqna9j1
+REl6StQ3LP8Mk9M1zHjNQim7eenPErRQjXgYE3SH1OqAiQZJHH5OxvgagvJ5lUl5CapZXFuFCo7
bPOnOi0PkI9n5UAhW+VehHkZCr0l9qIMYJ/Y3qqK5bUvJSpm0ngPFOs8uu0KKV/VYvAEaJSI9HDx
8rV/8rsXiw1vEpvV6/bTIn762qIGpUqTLT6BMFe3WdMDpkFPHpfEXwNAhvo0Lg/Fmzz1YcFfY/or
XzrtZL7+JXa7NLsx2QniKxs9Y+8qFgYoAx63nw6MrlVfts/s5BNSOqyd+ad7ib9O0DkW4DAypwK/
o6tRQutWbCC92mxvgmrloY8GtNUt+B1VuaLu7m3YnOL4zQIAoszDPVOY4kn3VSyZsclFg+DEPfag
agSBh8+i3cQ9nwlJjr+QsovM8w+zLPVQtmFhLepwmAglzyfCQVeqsE7kPybyxojxUc6bBvvDVEWn
4DJvnFpv5EMOiVNEizSPRYOiwkWnSJB68UvvmsxHb0wXbQ29Coam1VGmCAhk3wa/gVDF8sKw9geL
f+VCrwOkTOd1Q0ffCK6/MSBeuKIRAmHlktQX83Kn0RSwP+IkKYFBTE7J+59hvSS5d+ZZRBS4LwRq
dh1IwM2YNMQRAZobqr+sUgK2ZjmaT+kFbcd6/Ih1rS+Tq9nYK0IAqcWeglb5Z0BoimrY0ISgqKli
sAQ9cLTQQ95hfc3ZUP+iPkG9YhRHD/e+6310/tjxjMwV9QgQT+2Hpq9egsHhA+zGC5lgJ+iXc3dY
x0pW0WbDNIMuSi2AQutVOBk2tXlD6GNjLbrSHyJWzuAuWu+gOZ68MZ8su/l+xAYRt6rEzFbfX/hl
hP41JNhe5TXsgoXxDXIeG3qcZkGt90nhxtUP7f770PYASq8pYQUSk+TOPFpKYkH6Uy3ZWuO0HB/u
44enQHVmL5wQSrj/tjO51Yer86XTONNFIxh7BcL0MqpWIzhiMHcIxWt5NfgHB8jYSxJwKBS3SHWi
lXAQ2S0sVu5ldP/cMZsglHa0JdmgF5O9rWw13pYgLTtIFBCbanat1INdLRY5WQjOMR4uqBBQyHvY
UyNHLW8LRshcYMhNnHDb8L0epaAWQGYdWHOJVcPGH9oxmyYVROqfCWTwtAvAPbXSFKJJQcnbRcBG
12YGH1PnHFTdm3tHqzNodZOAMcD+Srz8/NLRUK51qG1GzfgPvWqZHG6Dgn8cJauMvJ6SsgK4QKO2
BJsH9ET41bbzYKbqcx3e1Kbax5pH6rgDspVYOn1hG35UNY14q0mg3f0yUEyhWqUUeIPUnBhQY/lM
j7aiuNUmqXDhOSt/ShruO1RjLYZtkCHVyck6J9uo9oh6NFDq56M7LwOGL1kYNpl0NF89rXKwwc20
CNjUEDgXPtuTLwxF1l22ty2dnllwg913VSzGf9mXBST+1MXIUpaLkbZvBmzUXwIgJuSMPdnapXi3
qZEwfwix4TQ00eYgqiuHWp8/05D7gKgA510wr4fgt10ZaRcddfg2jBmQDRhknsk3h/aoNUAGzXaL
V7RquFpVrqvSwyk8RrDjlTEaVlq23+gxrnL+e3xicgZXUK2R0E9nd5CuY/L7SQI1v7uZE4+vCsJX
cvb/asdCGqgsIWhxzleUSptC8O+WrhtbJ9W/bNFuC+U6ohFHoza3BkjvtybGysMda/HjYZOWGcDl
ipN85B3YbwsxTGUoRmVfBvGWaim0X1JbZhGbETt1MYwq9hKBB8cyRcM78APjG0+cybDcH+COZnWj
HBxteK/mDcWzvIx8RKsKINxQtNDUt3DlVrFqOB73wQ7VZx6Pu1Ht3wTxh7kO7nNmxjrnvbh1d0nC
1bZiOIQL659xUj4B10Vq0DOjTKEq4OEcfomwMRvko/zNK0MWUcD7M1w5iETvt9C3cBd+rTm9/Frh
E+7iEcBDdXIyM700HWQ/juDVOegvpgfCmyBll2HZ2wP6Rr91AcgcP4pi/pwTGbj8Y6S7x9aYsPQW
FDkn/FFqnsKUiQaZkHrmSEF8EaSTyykZ794DsqsCDqDuZi/E1c5yLs9IwLr4h92TfFVAmDBv+OEH
MlAIaZLjefURoBO7pG46z1DNbIlEDxqRGOrUJjk8klLW9JnhTKqgeTmx1tDVRIZOE6MhQboU9DZn
ajdlo4gyJL99mU/xmpf+3I/TCk/MrppXApPsmWn7s8ju4EcgMfePOWFVPfoDDUK3V+2mOwOTtRIa
Y7p2+NULsNqk5+nUfuFMYFdiV0a2ARPRAgTonJWUYi2HRUN5LsVlXdN/CVBEKfEs3yqNpsmjyBrF
oUiF7fXnrKBv3kb+iDdVtrb8K6ziW8qkKJNd6QjVkvcjrTYQu+xLMcHHOGdxksPxOTHpdO9qXIYK
X/4uyksWAGmItL+I7ANbGhyibNYhTPz45he2OLC66uwwj4+MOQJwQyzAu88paaNF8f1JXJDlSbDk
NjkdaEOk8qtVyQBhcsIcRy75TcHW82gf2dGYcj+CWq16Sj5jUEJTSsDXGnHPqRFTeIJ4/EbIq8nl
XILDKk1ORRR3ooZswce/OTr/0uBHryutE73aGsCCUtQqFll2iACEl64Oar+wNhc7Z3fXvAMR/eU0
65g2H3apv9M+ZSCl8kzJgUqPSBhqmDzfk3YDkWMBrzZRGg4FbH2fUtcyyT7KPRAXrpsnzFvJdR6p
FmSz4BA+ccfY7RofQpr4oOP1Hc59BlsVvhkuhWw1O3eLQ8KL6kLCzFI5R0jy7NM7a8UisLP/BI5W
bUrG4JdkDHGgS7JZrUfR3uyCpdIX7X3iJtI0B1v9yDJ3gjNorqLD7ecBtz4B/W/o2sYqLDJ4Pgk5
DHzUYUXO8KAalavyyr01S6D8ceE9ACpU6UPtFVMoxDlVAbKi4AY0ZZ1TCRg27kI+kqnzeXgKK68l
UekroEh2css0XkXCMVThd1JhGEl/tlXtGUfGYambYASVIodnGoDYm+8/QYL/EGZuhebPP5C1bYBw
tp0DNuyg+QQWZiDrSDmp4Lxj1xbbH5cw8BO3CsVj8HuHZiAndzlq3q9Rg+4ljMqpOVY6/4azm5hW
/sBWB5XupVI8D2aFfMQvkWexwKvpNIpYN2750ZA7LJmqw3YuhHDHihJf9LNvrYawj7xFxS/E3w2x
XvSj+/ayIlj3UQjS7cWmZQgZn42zR7/WCjzAGjqfBfghbB0fvZ16FH/BBSxeL6etgcsuOvN7ZCgN
UcxDQKsXFHaUEUY39y5vjGixA4QxRpUPSm7di6dnt7wv3d504AXkf+ndrr/IatIQ7clEAmrONiFu
8FEOTE8MS8uJGA2wRG3DzKlyQRoERUAXzx/ELJlJjeletwVKT04b2zMAKpG+0cmBp1AZY6uMNHMh
S/aWwwJPtMnemAiRRvjbq/BYrsZkMA7lwektH+j7GIdZhUSm+WuCOeYtJyyvvHYZTT1i2VjWnbuE
H5HzrmYI6YR/K16eGpQjzEAEyCIw5VHrsugzz06RLmMTnHZDms+ZtRCl+bNJm2KPT4x8trjUt7MY
D/fGGLHJRF0PSTIsWQPCGrTGKgd13uiVQmCC3mvkNVxe5IjTYeCuFx8jXjQGNQyQy1DCY3r/ucQx
ztXtsh9KChaQNOel8OGqyIksNg3rbhl3WMQT4uuF96gwl7nSN+I5O3rcne08hPTLxWwfzOX+r0wU
1lqK+kLxT4DcNNkAR+r2j7aDmm7CjcCHF2zgnz8wtw1sKKcmtH660pAGeM75nvIgHomty4m/vpJK
mMo1FQqQKIasfbAoVdW6JfMeuxo43poJKfbOBsfbSvw6bUbRUk2V71I9BMgBG8aUz0f2F4Dw4/5o
MPxNhxpg4ZaKz/qkDckSi855ZgfVYxSlVZYEo4CLGdsrZiuHJWnpWZR02n7HFy2INiFpPQ8HroUc
Bh5Bo1OF5/D6OgV14vEuZFqr/+uZzsD57j+krp1tB8Dh7QuDWknh08MF4aI2oNj2s61F/co5XLgY
EAZoRq5lNepEam94xdePXGiIxOXr7qWxcp9Qe4lrwvJwy/QHmfyRzJBdtVzgipgeMhT3SEKbiNfk
zzvuCDXGwoOsBlzZ92/rMEVG17/iN7GE0CxFYNP+QaXfALsxX97O7eORTblQxet6Lr9eRRZxOA1G
dIS2FzxS85khgL7U/1LwCCNh5srtUDx1P57bBb+P2r/L4lIalvJEBO2fcvY7vqoLAqN5cdcgj8Yp
IfIlqb5Cr+RWefTR+HCw/vrD9zvjG1SNk3eTXhOOaQfuUuyaPgX+QBBvGxmP6VDlYqzFp3LRzIXP
wxSsl/fpihNS2FBt8LXQPo+q40Cfr34LZOg4HS3Dz7GpeAgsniev40Xf6GOGtVrzNQq7e4LImK0d
AMh2wAC1UOmpGpnyuLgnEMCipzEtsYEAoSDU11wnj19iiz+EA93pfJg8G+1DRro8TPvrsUlRqEGd
g07gPSqJOvNy4KYDxQ7v0UcisNXxN1rJhI2L31UOFFjFtRSJ01TjnsOhaCbMvWb8+51nwtZL/6ay
xOkjw8OGpitLh8l4ZO9On2v470gUyuCX08HZKisJrP8JLtzm15ArphRo15bNLb2vRU+t7gMot+mj
pkXapR9cLSGgH+NlTPUAM/AKHVDe9yWLfD0pzZkaH2VwqVNx+l0xi2y3MMSAj9QlcUnvTrROS4FI
kBF7Tpqqt6+MX0bIlZrEccQdon0NT6nUAVs5Bt5uW3wLgL/ei2bBmvJpwTYAnnFz1Uqtb1CNKaYr
Q8TspucDbYpcYge2aLX/nFWiqBBZKlK5vVAHG9t5oduXWZ0ngiM/cSosE0zJ5eNI+dZeh8kC8RGn
n4YZ9yLxh0nJK4hAlSPg1moZmtLYcSAEwDv49bqXfSGeECI6ZUFJNQzvXFtPp3sZ09D9A2PVS16s
yDFtNFUwulp2GiMTiVHWZmNTydMvf199ls5aky9Yd53jEeiJ0w8O5cBv7YIWrTS5wGiwaNmIH2P+
zA4SG/4RVDTeV0r8CptO2BKupETiEKCZBPg8t8NvPob58QV5Pu9O9gtacq6t0TEbVY0/l/2DomYa
lHoKU0NaVf7uPkrAMXnuFBGIXhjgqDUp6zLLKkO48zBLkiKTZUsKH0Eafw+PSHU7JL0AfMuun04V
PKdLGNJK0qIuMVkcamXS53+Xq5eqL7+9GTMFIPtix0FwQbeVsd1UD6T/iWULtubdwKTZ4BMh/2Fe
s5d9Qnl22L+THggoVOrCipAePbPjeF8ihfTjzzWX12krN8leXV3bmzWqypWzbcvjOX2qSIaxTlze
eaWKutPYSWFfKRjBXRGyk/n7QbX+U2fXGqFUNzgwLY2I39/ofJNnmQEbstasxJWX3gMW0E2eWSdz
qdYoAYJ40c6aXr36KS9LleEEBWAjqGj3LgGUpqqsY4qIQd89kEN+rEuAy/icpfrlAc36A9XqEvxB
mTxHms8pzHkrnfz9DU4oWOdfAMzZ2Ctkf985C2VEnmSE9Xp0TYeS7iJAmmboGQAogqSjgbLAJSM1
Vu1LjYsAa09Fe6MnAh77zNjlw+adygzwxyFvxOT2JEjz83rKYrNgx/7vpWnPGKY5UkB5s/PBrPAS
IGYJdobCaWSJJgF3FCH43hRvkHvx08XDfyVybI0gp+1kQmyt9PgEXmSGPkI9CD0BBjda1w78RooN
hLa4aQfpU/dh/tWCNgBuELfBetkUuhjVFqJcAxKo+2Nc6PI8skpNui9ahzt9OMilJgFqqgPMS3Od
kztPlAB+p8r8CZ3kBXQ7RlN53RRfI0gllPjC8olrmEGWMvpNs7mweEGd1ZAjV/d+8iESh4j7HLNS
do9C1d7zthJy+bU+dJ/ybgrfXW/5qfaL4eSYNM3HU0h+B8/rRb1VY7ZSPGDKgO+qlkw+5u41hqaf
4PcyT7Bqj/0xH9QhTMOF5FPG1Foze6RPuPEQfMv4OvPaUaPn8mr/gE7ah2dTd4JorsbMv1AnNcw6
DYE0op2XvrXOiCEusDqWdEBYFEOd8x65nrZanl33+Vkr1QRoOE3pz6TskgAm3h6wLJlCRnWyGNdS
3xCKX4LrZEjpnEmDUKvjs1/A8PWVDRC/lfUA3A0jIj7boLPumsCXG7tXKGjBDB5Fz07Eo4VoNyoL
fa8jr8IysKcHMSibsKBHpMObKDh/ZN7Jh2AO5RzssoghMrRZatFbgWYbajwyEuEtTuUNgx/xVUhB
WuSHTj5RtDRgxhkkAximBR6zN/Bf0PGlelEd6kgErCl91dnOmoiDC/axMI/ZuZfnFhXcQHYcAuHU
t5PlOYPR7OaeYQ+LZ27pEEwCGWY0ARa9nUW5jFBwD7UHAmCswbcUTWFoz2vmVS0x0kDqNliUUduK
BW28gNnOwprhzxeW7RdDDo8Bm9AjCKKGoWb7RIp5iIke8K6Hjv7GXWupuLlmyQaOyHRQndlqR4Pc
2UO6FKJ+xi11F2D4dLTUOfAth3VOOr7y5GpIggYSN22C7nvFEuO1WqIWlodogLWUqJyTiKt6VFdg
l8EEE7TsvzmwxrF/6JrYqP+rPikVVEPQJNQdEidOdR7LFCyU4UQyVB18OvvNIhwcXnf6IwI3Qigu
PlxAd3uKE22JEp12w+dhsMbMKjrTgU4W2RtuBWlmuAt7jhuRPROLh8el/px6TBUS2ZxgV9CZiWPS
y6iKslBr9TFOFzx8gyIZ1BhpFZnW39K8tWPCQwLgkD1hUk53lB88cStaS+/mkhBCFcxAZoFB2W07
k5OzDptsnn4P4Zjgue85/I23B0PWCEK5kgo78Ir9bugWKusbklFcQVzVY629E5Ho5vmJ/m9mbrTt
lQbBMA+eMQ2wAit8J/Y1qJUveDncNb0BxQAmMaCtPYJJWL92c9d8JW8ZmRqRSnJc4wdwIiD/Tk9f
IPlN+7S/fy5y4TUlbWyXG7QCfBO0PnT5lOFiXwGCGIwjzzRZail6XyiXPUlF5nIKCp8Fx2bBer1l
No8aZJE1Z/zMwCUpbS3Im7usFHB8mke4tZ9XJ9tztYlLLsYznzvSR5f3/69T2QYzPRC7OwMxnUBS
x5QyEi9BJ25suAsz7Qtoe0PzzlJwb/o1Zr5OjAJbLLt/jDNL75KE7whZzHOdL64ygD2wzCxNkQ9K
jiZW9xlJ1qgl2u5swvLTP8eyXKpd3VIo5tj1qD9jreIzkJ0uAFS+oRtIukq3vtLZ+Y0P0Ts3az+e
UImpyhJcxhKCGNN3eAyzz+H4WrCqje6HqkSfShDZ+6k3k1JxoCyhnEl60w9y4gqPBXlrDoyc9DeM
e7HAx4PucqEoykqRns4nGjZG9biqENNluAXHXoYSaN/h2nHTCndN4JaKgXLr+kEFd1CT4ViL8mMh
sZpGE6z9gr3uOakSRlHv34lnvgMpod2gcazIt00UmE/fDW64cbLK2fm+7+j7AOyJi1hv4cocCzwA
/brTmP16h+AKT3a2AXQH7hRjmohE7tGyzVOpZqQeSXjumK5CvZqpv7DPjQLDnXp5vwLW5FfQteEU
ZrYh2vn2PDEPUEnFV1FJsTeeWpeXq+31DWPGF+eh3ULxwD/2VCkzf1dZ475yF55L7C12/5XLHnou
HqZ6exC6GIRPk6nLz/CSUq3yctywqWit/WQyiy9k1mETNv1QGC+2faxkxbgU4CWEeQwhZWcMQTNO
Oysn3b1ntH5uhxyXaMU+SZlI52Yy8k7FciAe5N3yBZJYD83EyEPStRe7vMYCgOh4XsRECTdOjAvL
dVe6Jx2/jP0XaVeNK75gaeko62JDvHT6x/kNwSxb6yLWMR+BJwvMPNLsrvUGzrqJaerrXUzk0Mj6
sQXs2qu+KOXlhn1PEQC4rdX60M1J0lTPYikXsKzEYGLgIluFZUG+g4jIbHCnb/HS7kSp3B7Cp2JC
sMHR0IVidkQVTMCJRm8Xz1+ihp2FY8usJ83AJfWGn/85pjVg+7PzDF1bDhuI3NtFJ3RSU7YNMgvV
ttYRCROQ3JaHAlCt4zii3+PrKW3EJr5Z6Zhsq9+3N8hsYXbEJEXVBJjVdTmMqAmsU46HwLnv4Kaj
bDT+niWcl+hwYFsY/oFY81wyxT13+dIGJB2Cw97SRWm2Ao4+1MoE6W7Df2bj2fuJpzi8exJ7kh0F
yKSADOF+l8o5n/m9EFlN+oD0RgWGV7jDINtAvDgsF6eFpyFH0mHT9LexC5NHPhkFF9VzSqGHER8K
ltM8hLG2WaDTWIiJKPguVVPB7YcbJiojCZsyCHv25VdSesl1ZYN1hTp5qdxV6OLr7TUFMCYgbmEQ
EawIHqXQdH2DASqT7dQXN9uxCIhB+S7IKogjiDbEK2G1mgdzox0xs3oEiWC1RSD1fCyTZCntBsYU
CZ/pW5LPsJ/dVh+USAPvOtFUuJJUjYkZpcBAlGcCSEVY42pqzKzr0NTJluJaz8m7L3f8Z5pKpQAr
IFToB8keJxtV6qQR3JEv4/tsYUItepfMqdwk/3P9INpvJBatNPakyC+7tYsPeWWJUsyIofpF5S3H
TcGB3VJAX9OggCfs1PwWEieL0+K4m0SJ7K/2q6ya/+pb8cEevuKUDBosvuR4iVkMMuVBVtWTFrWH
qGgQj9iG6YipW7l7Vo2MS28jEUSMLqamU2xcyoHqjUs85yj+5B+qg/lF+UQxojeG5HB9pndNtIEq
hCCyZhjXUZmHItQDbs/fkbkKW4RGG0cv1d3pYXB+E0Yc3mApX5Gcn2p+R5/3pDsjHE+fr0wCikZM
GdxDjUZg2eNV4Q0krRXJKH+ndsJOQ53q/NVcgRW1vlZM4FdcmQupKxq1oeUhRSgIxHxNU9VupSx2
oSYEsHQf/6U1Nai1syg/472gfoDn8GSwzLnUhAGlX9tkkqVW6MB5ts1wWNTvaU+xvTRF+je+ij7j
ficL3WaQqlmQ6BNp0uvDbiE1tNxsYY4n/ulLmESuFibtsqGvxFVEswzSY/gJHX5w2Stm4/7iLXGy
gKWkxCV+01ewpSf7NFW+k//y/Hzn9jMTxISWG56PARrK675q9/ElliadzBt+xNvry4NAGThf+yDY
AqDj4pkoDYoyNXa/0mqRm3iHoTapyvxohc1py34wn/LuNm7MMfKQg4U4hVvsa6iXyxtM5MAI++Co
gMwv3guM8dO37lL13PtpEZI1s0fNu26/5jcUEQ5Ei7DeeUfjSA7QDvJV0iBiwC/BKAuoG/CvOcND
pNX7+4AH9+kSKJs11+m0jAYLZLbtX4f7L2/LD4PriMJ0/E5qmvCSs8sWahDs3vw52P9YT1FRMOxD
AREyHZ5H/mSQNq4wsu3MuhQsiLZDZGnT8RQJN9HUHBULr7nHZ0rRaYWVhVVn90TvSi5t/kTQioom
yzleyfvyakahx1b257o/JO+eMxPXxoWnlnRlAaIWcJcy92UJ50ZW3mBf3wp6bguOVef+OS7DQ/Cj
bMSaetB2hmEObepNp2i6hDV5MI79KhNa6OdyTLQMBd4tL5NeibQsxqlK7N1R+YAkZR7nW2y3LzE1
BQhtbK1hmab/UkW5gjU9e9OrFKjN0A5Y68CyG1hz7rAyty8L6dmZUndjuusIAWRgVTmBQrypaY67
UEoEzRXmg1mCZKWTkZdzjlYAc10XkAtojB/zB6dci31D0l80P29tIKWAGgQ8bTn1gtEQ64VsOH9r
a5EAvKEFhmsYptGCMJxMQaCCDeX9WRDHOZeeHSAb4P6cjysE5rw1Mjp/kvDqnjOn09VxUGPBnLjR
wopyz3E2J6+4VOidDiNKHsaHDxv+UIUvXoYBPjHad4e3EsW37HSt0CMW4s3LogSiIasRWyAYX/cx
72rVNv/4uQEkcufPqIRjyPGFaDCD5xAu/TQYtq6xP2UUmjJVh85ZnpNk7rW1z7IxLIBm6mwcbxOO
hR1FHfCl1UPYEC9DwS+g/sZGuyDRTbnBdDZRP537Yi2edfvvVwLxR+lJUgFB0gLVOTWZZ9uzJBht
PPygw2c3Uc0aECEisvN0oGKD2RCsWfKZPhuyOxnnHxnYd2Sxhyuk+kWDfT8Ss7E4HmJPWV2OhKsX
uKo6t/EcJ+l3pC8pIp4AUMryot5mUOoasBUaTBKoETtLweT3WpnmS7+sh+1xmL4THsHZmL/+vBzu
TvjbpAcerZvJoBHeO3x2LcFp8FuVo2grrMs9Mz0yH3AiwjGO44FXzOKSP8+R44daW7ezQHbqi1g3
VutDlWaRtm0CGWormMLcz+hVwg+4L4XaJSSiRFsRSO3EBi7ok/Jv1MvKYXJHgf5d6U5ASk/3f/KS
rrKC5zzC9xz0aW6ng9hhjGG4ghDWDTf6VI8hf1o7u/O04ogqEkHggxfUq7sP1fJMl6dcAsy78JTH
xvuLwb/mnEHjL6tyKEIkuf77pcUM+62i5/DyDho8Pu126HZRLpFnAKLLyvx1ngkoeVdenFlQddQx
aoFwWX2MVT+x8IIPU77NHeplqzDAD1sEDBgdVbKc3FmIcIwa1lhTmyRAC6NXCZHBGdpAqjQxOf+g
przC66yugiZNdO2JkDwwDyr8jEIduELhIIV8eanWhdFdmergBrvNhb6Y9KAPuv2MyDo+1tA2XPzu
80HTumSYcLLm/qN0Vl5iRQq12fwlDemj/JAocNGit8PwPwjSI/4/UgSq1LMt/7eQu8bDFwEl9SLE
mmmgzGb8gSEoBM++f/D9W6e8a0GUplNNS18FcOGcJSID0kmJs7EBW/ZTfsqUDOe66k8RaSJ8cWiw
xDxwfweGceStkYtl0VpLZERzxSO2aGStin1WNtYiU0aL2q07+1BONiGtveA3D+VuK0Rxeh8pjXpl
TSJs5LsIS63LWUXkdv2QpA/2QjN1BCFbYrRzAp9BdByBmjHbzSy8KDf2mPH58I04WuzQmsukJVw2
54KmdzqAIHqv2KYPv3mJQ5cb0RwmeDsGrk5RpRwzxyzX5DWFC1QsZzt21dbf0xK4Q9QzwIRg4f0V
+jEAmuyCl0og1uKg1zKkho7qyqVrn0QkCNV3J4OX0wENdouptB/kf3mXyvpjJ+IwcYUZbvmIz746
0VMzmGqdaIAbyQGTRHksyIpuhvVNrX0Z+GMdtWIYBNl6ZNDdhfJaA29StJbsLOtfxpMB8nwbb8tt
7MOuX6fG1OZL2RzEDS+R10JhwQWM7ST/l0oHaSj4YiKJV4gHlQ3PP4Jw8WQwvCE7rLQnyBREmytK
RPob1eW1hXOp5kYBJME/+D8SCnO0j7M0lvDjSya6VuxnwQzqzL4BodvjYJHRhNcrN0DdDlYj1uSl
4roz37ym74tOWrEKnWpHlsrzRAYWnDTf7iGfAbhv3zy+EpQh8lYc+pZ4OU1NO1wMvCFXwuTy6Ves
eKLKKys+fGb3J6MmI/c+nIWR4eIFDmQgPtsMyjCgzF7uPsGHRmHmYiBLVuMaDWX5uVEmWCEyU5Sx
QS4OTGm/PdBoTRw7Eznv9RQAewLYLC1vuUzHfAzqZnI4eJt4t4AM+vRtixg63xgymQXAmPECXB4/
+YKElPLXSUx9e/p1V2OX4fxsuKj6gCBpKl7WpPWDHaejHlx6k2y4O/KCvCW1ukCq9opezIzRQM1b
MCO1ep7KwZPfji3JsYkDX4RznmPuzqxeOah7ROPkYHdd2WVrV3FPMZhbNugThHxG+mgWW7DZaA1d
8YOGIm0+6iXVQFZBoGUTRtAwM61uK0LX+qTI0Emxpoug+8rcODidkzOGFLcAzxi2Ln2cL4ezuRnq
dRyiwfFUYoiRlIHyqUrggszo0vnY9784lK1zl1RVvcCXfT4ddSwUZQ8qHa5MvjfV7H5jFSU44rDm
qL73yfIut/E4PxAmAUdYOIDQwPu4wxJHyW1D/6pMSU0J5Nv3NIj+0sukLiIpISRBVCe63HMUTL+9
Hr2JGdVTmxg057+SyYgv7vA3u5RFCsnnXpfLbyu90iL9+CkuTJVkI+Y6Tu3EwrGS35GuZ223FKV6
/loypzxxStPiNLpDHcxSKLjtJKxu62Es37nV/DvJWYzmryDMogBn7afhU6Rlwp//ruwWlRL6TU85
HE5Rbll7N9ynCHUzRLqHbUKjdS8+L3FmYwYqgwf2alwCEjxEvGus4fTis0W31t5xTBKWsn32uoJO
hSRRACH/mMA/LgCrinfMFxqSGvm1shSKn9s5qaG2pCr+YvociN9/xgc6JKz+kRj7J14RB5pSVGlZ
96fcUBm+gHlWyU5aRO8jgYnBcgcZV6vtsWTeEi9vO+tZdLqwdV7LeQIWLW1JIp8JSpmb4rhSrnTw
g0N6/nflc0hyqfMbtSdSm4dPYVMbyWRIvGfTM3Ay3VXMv2eLzDOVzcQjQ5f6KE9BE69J2gv3ayxY
t3sd7qwcC+64LXK/zIl7XCILqG89eqtOWflwxWQPxW6vKZqCJrjntL+UuqajK5W7XJ+Rn4GZGxlz
fN1nljgv9vRH6Fkvy96pSlvhVediEFEwv8e9zrgMbqIAUqKgrKHOzY5irdpG7pLL3rldAjl+FF9N
J0VA3RSlh9BTtUsFyZqBvR2bYhRflppBFAsVHdKQiN6E3zbhypHQKo4INTDipFpjT4D4hHnVlZU6
uIM7G7VP0Vr2yohi7KsmhnUscpUoGRo+V6H5Rras8aYzbQX+Qt+IUTAu6CflurYztziC1AD23+C2
CM78FLKYeWhakIlP4v4U0Y/Knz3oVOg+4EHRadOAmhjcd56luDCfxT+vdBUELv562kSm7/G4Sqyr
gNXLldeXjwEtynxenclEV+kDs8yasm+p4xtSsnpOp0bAA8s7/LTkjR0sKa8k5ohELlg3UORDytU4
J7c2RN7+C6hvNAM2e80yYf/x1vRK0HuixTe1wHigEd5vsvUWQ0F+/Fl4laimuBIB+bzlhmWJPpHQ
3MIcNCHnA30McLcmODnPPf65NWWcTNgj/SGmuRrXpfJNHBtLQjGDO/TPPx4uJf1hiJYccZBCkG/b
O0DBvdZQx3+tkB7+M/tUW23BrfUcNVk5tghnyfK5ns8p6XrvUOU1RSYdkACucC22QUq6NZxQA63M
kvohgciAyEf77V2V9I0pKHuOo2rFPw1lNPoT5zybxqSD93baL9fbN6Vwdy8PpDzVq/FQfbOXBIVG
il9yeJy8uNxLUVZsu1MBxdj3Ifx76J2fGJswWdtAavyss+rjcfB02fkoQCWJ73O7io8MyN+ue0H2
UM1rSXU6yYMT9X8iMVgXHcPtpjzNtNZ0GZt1ie8UA4WLwZgWMVkNoCjH30PjiACMfWHVgzRmjieo
kbPddZDIibm8O/tmHNZHbwxb9+bD8ht3HrlDhyW95o9J9ZNslTFJiy2pii3phiyyPr6dpPz8wOin
TydtpFN1zDdc1Ty1E06aoIizdIAIadrlJipL17tlZjn9/fDS8wgatjShrxz9aqLdWpq+G5PEK/SM
phmAJ4fI7D3zuQqEe3kJgQz0MqI1Fl+uoY03pSZPravZDr3CgR0o0ym4hDTxYewaN2Xy3QrNNdXv
qI9ZkZtwTagYWDAP4I8SEA/+C8V3CcWpO/r9wIWvtEpXbcRo9iA+3djj9fQQEIpKSCbBPee1jomY
DJEdDaRyNR/udL3qsAyyR3K17c57P+0mHxXxCykOix+t8PGKORD2DQ4il5nCPd7uMLJ5I6OcQn8v
ppKwNfnueuReOspitFBT1Hmb8aTgY2BqHsKO+wOCkzhH3azqlld1DpBvHo+wx0VWcc1bmUCJ/aiy
2+zqDu1UBNluZo4EtMqQ4DSCbvumpZaJ7GujSkSAH72CkY1AvOqb/3hN9coKqa5gcA7MKZQcDETl
j+5x4cW7CcS8XhJHkCJOv5zNmjE2OIlUeK+9Jj4vK9eiiAGjkkUEpqAMEsBDqXDhuboJgVywim4E
7zuFYrD0ZtlKUp7CI+vR4i3waa+FaYoWzs5cW/N89See5B7TItHt22a/Aqb5WX8gQAuLhqV0/NXq
S1LdDL/WoW7aPEM8IZuCKoyG7OPdLtYH2Di6LanAqQnwEeEOkVOGcUmcOvkXsCucEX1fQOC2woah
kYDY1MP3nFfRiwZcVNMlHHho9xX4+ZLLbQsczWG359862t9PQ7vlMWncHmVgcQYaaM97RNaNHIJP
JHipFBApnryhpxTiPr6nOBnRX0lhs9PdXXP7gluroJPkJwZwHmSmzyJ3sLyHUBdpcXKr3pcLuldp
jUyWg1/NY/d+ktePrQN+KjWrZX0fyZYVHpjKU4V4wYqMFt9VebaHlBIHjJgZAGWKv6B3POTeSvkE
C62u9On/+XE+bMwJ73YmbKJMl5X6+1thQXGu6JbQzMrT3Iq95k3S164zDr4IwnQmxkWeiCsx58fQ
RBVF9w89WthMAxNbByPFAfBIgRF2j+EOnXmebN/3QZC8ZzvIUwKAjejh6VEXXnR97+rFRQ10kASF
Nbdq1BeZmZwDJG2TJyYieubDfdGbkS5lrEX+FWZtlZyjeYud56P3U28ybwvaJsFJt34e1AG81mPk
XfkaLt8Jx22sqB9Ucp5Y+P8wqYLWMolcp7Or9HiEEm0wZZtRoUSsEaWqUQ6v3U2ZaX73Lxh9Ua4F
kWlmxIRWegEyxH1BYPZ/SjA72p9hmGj4muycsFxSATaPm5+eBy9PNp2TRozmJyNjo0ZlYpvULLwK
3YvJ6jZXKwB5PBS6R64hzCMioxnFlW+73eYSSnmsaClbgc+H9dGWcjzc2WsylmJ2vPnMbQyv0FFo
A6ulkQdq7kuP4vOAIgXO1sv+UKe9RuAs9hTExr336rzMyIyeK/BQ18TO6H2i7RaffGqyV4NM8psS
27LRLlkF7kliqQ7XbHMm691dEYx1KslwHxkaLDTzrtrqEeb9Rl1GKWjCa85sq+2uOUzFcscfTUaC
2iWgmq3hWz2B5c4KMVxKizPaHO0njjTHuVTAG8mjuL5YzE3Do6X+ZpN/3JrH5hpcMnx/fA7g9D4D
loWpiCJM55tYLho/R0ZgJr6UhwyLx8Qkyl9DUBiKQKdqHOtB/6LfJxoxZ40ahacgQg7gOrvHOQXw
JjJFbvXIS974s5nWAQ3l/vQ4jEgp5aiX95fJK53cSwcayvrBYa5dpljegxdRLXayINhg7TMpuIB2
6xyMVnmVLOowrRL8c7mbZZIDMcxkyygIGldY/G4ScOWMhO0jam6zyCxjLg9VFPODUtIS9JJfBjc9
lH2Qwh4YMllY2eDVf5vvrJ7huF8iVCIFD+h84yxgb7sR3+CYtTWMlQL2tMxc2eIPwkJY/vvSa/7W
2jRQS1iMMFBFBe3E7nxeHo88M0JL7RaDOrs3QPwJ/r2YWu0w78YSjR2ke/pauOT6C+P5c6KaXUEF
fGIfz1r6r/pteQN4/BGl2ZpPDZ1t3brUOT2rPljmftqtni/IjB2ywBcd6erWgzCygKfUfdn4i//R
ysEGdvMgLNgYSqmF6znK4TroZmokX6Ls5al/Mh0XqqEcAAuep+z15L1rAWcVYkDjUn8az9dKvLjS
AlKkmEsd+RZI+WeWgqOoCzJo76eODJBtpSw8theOqpSBLctN0pRtckrafeKMtQViZDzBDUCMQGeS
oQMfoT6BVe5BJBrVSS+edFZPHgYgZMyS+AbTFan5N7Mok6XAphanuPeFtjvvtOD9vtvt9sdvEDBR
3t9niAlkG8LtQRU3H9pl4nL1imb+L3osVT4J7CT8L2vnNI3wbwW2qeeX3tdcLzS3t1p/82nFTkol
7q6siTPeMm+vdTMNRCn1UqXMG6mCB9ijwnufWpStLpT9v0n6xf+d2+Q1gT2MAZkW5R74OPDWAJMw
tzEl3TCaQohLicApbCYHcuq51t64jBm+yEdJVjmvJEXtWlzB/qP3PgJhPbfyJBFL/HRMEoCi0ZWe
IUH6vS7GmCRua155UeNngY9Fg1e9oOfVapfiMFbUDq2NPU1GydsV/G+ZWXzM2NqpwOOIPYB5cxOo
h3Qo7ctRUkb7lOyn7GbwuTcaLz1+pGzPciB+SlYwWf5rfxBG6m2Kyb59pe2h19p7MhLb+xn76DJm
0lTe/fvkUW/hdtQirxhPOhgp/gtTyTLfsTEiks2nZZ68W1pEgtutFyDz7t/yfAPXF7cRgNEYX/ZN
Ze1zmnU/20B6vjKpBFmCOKRlxoGZTVCTk2kIRqBRl1OU6ieo/mjgbG52I0MCZp9oDf3YIZ42BeCs
/3Ae4a0VaGo1CaCCBA0imsqhiNBmKbYNACwmVDutwX5eWoR8MXybc0is29g2vmEqCj2bkCwNWz+t
KOPouE4CjWLmnTqnr7f3/8RNtVTDkqKsFJ7JvTAeaySIKMuz/EMNQuqssWpzmDDCjOVWXtKXaZNy
UYcMA49NisN6VoKlKHJ9Og==
`protect end_protected
